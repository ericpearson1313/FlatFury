-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_enhanced_pcie.vhd
--
-- Description:     VHDL top-level wrapper for Verilog wrapper of the
--                  axi_pcie_enhanced_core_top.v file 
--                   
-- Comments:
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_enhanced_pcie.vhd
--                 enhanced_core_top_wrap.v
--                    axi_pcie_enhanced_core_top.v
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.conv_std_logic_vector;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------


entity axi_enhanced_pcie is
   generic(
      C_DATA_WIDTH                                               : integer:= 64;
      STRB_WIDTH                                                 : integer:= 8;
      BAR0_U                                                     : std_logic_vector(15 downto 0):= x"ffff";
      BAR0_L                                                     : std_logic_vector(15 downto 0):= x"ffff";        
      BAR1_U                                                     : std_logic_vector(15 downto 0):= x"ffff";
      BAR1_L                                                     : std_logic_vector(15 downto 0):= x"ffff";        
      BAR2_U                                                     : std_logic_vector(15 downto 0):= x"ffff";
      BAR2_L                                                     : std_logic_vector(15 downto 0):= x"ffff";        
      BAR3_U                                                     : std_logic_vector(15 downto 0):= x"ffff";
      BAR3_L                                                     : std_logic_vector(15 downto 0):= x"ffff";        
      BAR4_U                                                     : std_logic_vector(15 downto 0):= x"ffff";
      BAR4_L                                                     : std_logic_vector(15 downto 0):= x"ffff";        
      BAR5_U                                                     : std_logic_vector(15 downto 0):= x"ffff";
      BAR5_L                                                     : std_logic_vector(15 downto 0):= x"ffff"; 

      CARDBUS_CIS_POINTER                                        : integer:= conv_integer(x"00000000");
      CLASS_CODE                                                 : integer:= conv_integer(x"060000");
      CMD_INTX_IMPLEMENTED                                       : string:= "TRUE";
      CPL_TIMEOUT_DISABLE_SUPPORTED                              : string:= "FALSE";
      CPL_TIMEOUT_RANGES_SUPPORTED                               : integer:= conv_integer(x"0");-- 2

      DEV_CAP_EXT_TAG_SUPPORTED                                  : string:= "TRUE";
      DEV_CAP_MAX_PAYLOAD_SUPPORTED                              : integer:= 2;
      DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT                          : integer:= 1;
      DEVICE_ID                                                  : integer:= conv_integer(x"6011");

      DISABLE_LANE_REVERSAL                                      : string:= "FALSE";
      DISABLE_SCRAMBLING                                         : string:= "FALSE";
      DSN_BASE_PTR                                               : integer:= conv_integer(x"000");
      DSN_CAP_NEXTPTR                                            : integer:= conv_integer(x"000");
      DSN_CAP_ON                                                 : string:= "FALSE";

      ENABLE_MSG_ROUTE                                           : integer:= conv_integer(x"200");
      ENABLE_RX_TD_ECRC_TRIM                                     : string:= "TRUE";
      EXPANSION_ROM_U                                            : integer:= conv_integer(x"ffff");
      EXPANSION_ROM_L                                            : integer:= conv_integer(x"f001");
      EXT_CFG_CAP_PTR                                            : integer:= conv_integer(x"3f");
      EXT_CFG_XP_CAP_PTR                                         : integer:= conv_integer(x"3ff");
      HEADER_TYPE                                                : integer:= conv_integer(x"00");
      INTERRUPT_PIN                                              : integer:= conv_integer(x"00");

      LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP                     : string:= "FALSE";
      LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP                   : string:= "FALSE";
      LINK_CAP_MAX_LINK_SPEED                                    : integer:= conv_integer(x"1");
      LINK_CAP_MAX_LINK_WIDTH                                    : integer:= conv_integer(x"01");
      LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE                       : string:= "FALSE";

      LINK_CONTROL_RCB                                           : integer:= 0;
      LINK_CTRL2_DEEMPHASIS                                      : string:= "FALSE";
      LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE                     : string:= "FALSE";
      LINK_CTRL2_TARGET_LINK_SPEED                               : integer:= conv_integer(x"1");
      LINK_STATUS_SLOT_CLOCK_CONFIG                              : string:= "TRUE";

      LL_ACK_TIMEOUT                                             : integer:= conv_integer(x"0000");
      LL_ACK_TIMEOUT_EN                                          : string:= "FALSE";
      LL_ACK_TIMEOUT_FUNC                                        : integer:= 0;
      LL_REPLAY_TIMEOUT                                          : integer:= conv_integer(x"0026");
      LL_REPLAY_TIMEOUT_EN                                       : string:= "TRUE";
      LL_REPLAY_TIMEOUT_FUNC                                     : integer:= 1;

      LTSSM_MAX_LINK_WIDTH                                       : integer:= conv_integer(x"1");
      MSI_DECODE_ENABLE                                          : string:= "TRUE";
      MSI_CAP_MULTIMSGCAP                                        : integer:= 0;
      MSI_CAP_MULTIMSG_EXTENSION                                 : integer:= 0;
      MSI_CAP_ON                                                 : string:= "TRUE";
      MSI_CAP_PER_VECTOR_MASKING_CAPABLE                         : string:= "TRUE";
      MSI_CAP_64_BIT_ADDR_CAPABLE                                : string:= "TRUE";

      MSIX_CAP_ON                                                : string:= "FALSE";
      MSIX_CAP_PBA_BIR                                           : integer:= 0;
      MSIX_CAP_PBA_OFFSET                                        : integer:= conv_integer(x"00000050");
      MSIX_CAP_TABLE_BIR                                         : integer:= 0;
      MSIX_CAP_TABLE_OFFSET                                      : integer:= conv_integer(x"00000040");
      MSIX_CAP_TABLE_SIZE                                        : integer:= conv_integer(x"000");

      PCIE_CAP_DEVICE_PORT_TYPE                                  : integer:= conv_integer(x"0");
      PCIE_CAP_INT_MSG_NUM                                       : integer:= conv_integer(x"00");
      PCIE_CAP_NEXTPTR                                           : integer:= conv_integer(x"00");
      PCIE_DRP_ENABLE                                            : string:= "FALSE";
      PIPE_PIPELINE_STAGES                                       : integer:= 0;  -- 0 - 0 stages, 1 - 1 stage, 2 - 2 stages

      PM_CAP_DSI                                                 : string:= "TRUE";
      PM_CAP_D1SUPPORT                                           : string:= "FALSE";
      PM_CAP_D2SUPPORT                                           : string:= "FALSE";
      PM_CAP_NEXTPTR                                             : integer:= conv_integer(x"48");
      PM_CAP_PMESUPPORT                                          : integer:= conv_integer(x"00");
      PM_CSR_NOSOFTRST                                           : string:= "FALSE";

      PM_DATA_SCALE0                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE1                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE2                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE3                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE4                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE5                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE6                                             : integer:= conv_integer(x"0");
      PM_DATA_SCALE7                                             : integer:= conv_integer(x"0");

      PM_DATA0                                                   : integer:= conv_integer(x"00");
      PM_DATA1                                                   : integer:= conv_integer(x"00");
      PM_DATA2                                                   : integer:= conv_integer(x"00");
      PM_DATA3                                                   : integer:= conv_integer(x"00");
      PM_DATA4                                                   : integer:= conv_integer(x"00");
      PM_DATA5                                                   : integer:= conv_integer(x"00");
      PM_DATA6                                                   : integer:= conv_integer(x"00");
      PM_DATA7                                                   : integer:= conv_integer(x"00");

      REF_CLK_FREQ                                               : integer:= 0;  -- 0 - 100 MHz, 1 - 125 MHz, 2 - 250 MHz
      REVISION_ID                                                : integer:= conv_integer(x"00");
      ROOT_CAP_CRS_SW_VISIBILITY                                 : string:= "FALSE";
      SPARE_BIT0                                                 : integer:= 0;
      SUBSYSTEM_ID                                               : integer:= conv_integer(x"0007");
      SUBSYSTEM_VENDOR_ID                                        : integer:= conv_integer(x"10ee");

      SLOT_CAP_ATT_BUTTON_PRESENT                                : string:= "FALSE";
      SLOT_CAP_ATT_INDICATOR_PRESENT                             : string:= "FALSE";
      SLOT_CAP_ELEC_INTERLOCK_PRESENT                            : string:= "FALSE";
      SLOT_CAP_HOTPLUG_CAPABLE                                   : string:= "FALSE";
      SLOT_CAP_HOTPLUG_SURPRISE                                  : string:= "FALSE";
      SLOT_CAP_MRL_SENSOR_PRESENT                                : string:= "FALSE";
      SLOT_CAP_NO_CMD_COMPLETED_SUPPORT                          : string:= "FALSE";
      SLOT_CAP_PHYSICAL_SLOT_NUM                                 : integer:= conv_integer(x"0000");
      SLOT_CAP_POWER_CONTROLLER_PRESENT                          : string:= "FALSE";
      SLOT_CAP_POWER_INDICATOR_PRESENT                           : string:= "FALSE";
      SLOT_CAP_SLOT_POWER_LIMIT_SCALE                            : integer:= 0;
      SLOT_CAP_SLOT_POWER_LIMIT_VALUE                            : integer:= conv_integer(x"00");

      TL_RX_RAM_RADDR_LATENCY                                    : integer:= 0;
      TL_RX_RAM_RDATA_LATENCY                                    : integer:= 2;
      TL_RX_RAM_WRITE_LATENCY                                    : integer:= 0;
      TL_TX_RAM_RADDR_LATENCY                                    : integer:= 0;
      TL_TX_RAM_RDATA_LATENCY                                    : integer:= 2;
      TL_TX_RAM_WRITE_LATENCY                                    : integer:= 0;

      UPCONFIG_CAPABLE                                           : string:= "TRUE";
      UPSTREAM_FACING                                            : STRING:= "FALSE";
      USER_CLK_FREQ                                              : integer:= 1;--3
      VC_BASE_PTR                                                : integer:= conv_integer(x"10C");
      VC_CAP_NEXTPTR                                             : integer:= conv_integer(x"000");
      VC_CAP_ON                                                  : string:= "FALSE";
      VC_CAP_REJECT_SNOOP_TRANSACTIONS                           : string:= "FALSE";

      VC0_CPL_INFINITE                                           : string:= "TRUE";
      VC0_RX_RAM_LIMIT                                           : integer:= conv_integer(x"01ff");
      VC0_TOTAL_CREDITS_CD                                       : integer:= 77;
      VC0_TOTAL_CREDITS_CH                                       : integer:= 36;
      VC0_TOTAL_CREDITS_NPH                                      : integer:= 12;
      VC0_TOTAL_CREDITS_PD                                       : integer:= 77;
      VC0_TOTAL_CREDITS_PH                                       : integer:= 32;
      VC0_TX_LASTPACKET                                          : integer:= 13;

      VENDOR_ID                                                  : integer:= conv_integer(x"10ee");
      VSEC_BASE_PTR                                              : integer:= conv_integer(x"160");
      VSEC_CAP_NEXTPTR                                           : integer:= conv_integer(x"000");
      VSEC_CAP_ON                                                : string:= "FALSE";

      ALLOW_X8_GEN2                                              : string:= "FALSE";
      AER_BASE_PTR                                               : integer:= conv_integer(x"128");
      AER_CAP_ECRC_CHECK_CAPABLE                                 : string:= "FALSE";
      AER_CAP_ECRC_GEN_CAPABLE                                   : string:= "FALSE";
      AER_CAP_ID                                                 : integer:= conv_integer(x"0001");
      AER_CAP_INT_MSG_NUM_MSI                                    : integer:= conv_integer(x"0a");
      AER_CAP_INT_MSG_NUM_MSIX                                   : integer:= conv_integer(x"15");
      AER_CAP_NEXTPTR                                            : integer:= conv_integer(x"160");
      AER_CAP_ON                                                 : string:= "FALSE";
      AER_CAP_PERMIT_ROOTERR_UPDATE                              : string:= "TRUE";
      AER_CAP_VERSION                                            : integer:= conv_integer(x"1");

      CAPABILITIES_PTR                                           : integer:= conv_integer(x"40");
      CRM_MODULE_RSTS                                            : integer:= conv_integer(x"00");
      DEV_CAP_ENDPOINT_L0S_LATENCY                               : integer:= 0;
      DEV_CAP_ENDPOINT_L1_LATENCY                                : integer:= 0;
      DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE                       : string:= "FALSE";
      DEV_CAP_ROLE_BASED_ERROR                                   : string:= "TRUE";
      DEV_CAP_RSVD_14_12                                         : integer:= 0;
      DEV_CAP_RSVD_17_16                                         : integer:= 0;
      DEV_CAP_RSVD_31_29                                         : integer:= 0;
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE                        : string:= "TRUE";
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE                        : string:= "TRUE";
      DEV_CONTROL_AUX_POWER_SUPPORTED                            : string:= "FALSE";

      DISABLE_ASPM_L1_TIMER                                      : string:= "FALSE";
      DISABLE_BAR_FILTERING                                      : string:= "FALSE";
      DISABLE_ID_CHECK                                           : string:= "FALSE";
      DISABLE_RX_TC_FILTER                                       : string:= "FALSE";
      DNSTREAM_LINK_NUM                                          : integer:= conv_integer(x"00");

      DS_PORT_HOT_RST                                            : string:= "FALSE";  -- FALSE - for ROOT PORT(default), TRUE - for DOWNSTREAM PORT 
      DSN_CAP_ID                                                 : integer:= conv_integer(x"0000");
      DSN_CAP_VERSION                                            : integer:= conv_integer(x"1");
      ENTER_RVRY_EI_L0                                           : string:= "TRUE";
      INFER_EI                                                   : integer:= conv_integer(x"00");
      IS_SWITCH                                                  : string:= "FALSE";

      LAST_CONFIG_DWORD                                          : integer:= conv_integer(x"042");
      LINK_CAP_ASPM_SUPPORT                                      : integer:= 1;
      LINK_CAP_CLOCK_POWER_MANAGEMENT                            : string:= "FALSE";
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1                      : integer:= 7;
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2                      : integer:= 7;
      LINK_CAP_L0S_EXIT_LATENCY_GEN1                             : integer:= 7;
      LINK_CAP_L0S_EXIT_LATENCY_GEN2                             : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1                       : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2                       : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_GEN1                              : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_GEN2                              : integer:= 7;
      LINK_CAP_RSVD_23_22                                        : integer:= 0;

      MSI_BASE_PTR                                               : integer:= conv_integer(x"48");
      MSI_CAP_ID                                                 : integer:= conv_integer(x"05");
      MSI_CAP_NEXTPTR                                            : integer:= conv_integer(x"60");
      MSIX_BASE_PTR                                              : integer:= conv_integer(x"9c");
      MSIX_CAP_ID                                                : integer:= conv_integer(x"11");
      MSIX_CAP_NEXTPTR                                           : integer:= conv_integer(x"00");
      N_FTS_COMCLK_GEN1                                          : integer:= 255;
      N_FTS_COMCLK_GEN2                                          : integer:= 254;
      N_FTS_GEN1                                                 : integer:= 255;
      N_FTS_GEN2                                                 : integer:= 255;

      PCIE_BASE_PTR                                              : integer:= conv_integer(x"60");
      PCIE_CAP_CAPABILITY_ID                                     : integer:= conv_integer(x"10");
      PCIE_CAP_CAPABILITY_VERSION                                : integer:= conv_integer(x"2");
      PCIE_CAP_ON                                                : string:= "TRUE";
      PCIE_CAP_RSVD_15_14                                        : integer:= 0;
      PCIE_CAP_SLOT_IMPLEMENTED                                  : string:= "FALSE";
      PCIE_REVISION                                              : integer:= 2;
      PGL0_LANE                                                  : integer:= 0;
      PGL1_LANE                                                  : integer:= 1;
      PGL2_LANE                                                  : integer:= 2;
      PGL3_LANE                                                  : integer:= 3;
      PGL4_LANE                                                  : integer:= 4;
      PGL5_LANE                                                  : integer:= 5;
      PGL6_LANE                                                  : integer:= 6;
      PGL7_LANE                                                  : integer:= 7;
      PL_AUTO_CONFIG                                             : integer:= 1;
      PL_FAST_TRAIN                                              : string:= "FALSE";
      PCIE_EXT_CLK                                               : string:= "TRUE";
      PCIE_EXT_GT_COMMON : string:= "FALSE";
      EXT_CH_GT_DRP : string:= "FALSE";
     
TX_MARGIN_FULL_0  :integer:= conv_integer (x"4F");
TX_MARGIN_FULL_1  :integer:= conv_integer (x"4e");
TX_MARGIN_FULL_2  :integer:= conv_integer (x"4d");
TX_MARGIN_FULL_3  :integer:= conv_integer (x"4c");
TX_MARGIN_FULL_4  :integer:= conv_integer (x"43");
TX_MARGIN_LOW_0   :integer:= conv_integer (x"45");
TX_MARGIN_LOW_1   :integer:= conv_integer (x"46");
TX_MARGIN_LOW_2   :integer:= conv_integer (x"43");
TX_MARGIN_LOW_3   :integer:= conv_integer (x"42");
TX_MARGIN_LOW_4   :integer:=conv_integer  (x"40");

      PM_BASE_PTR                                                : integer:= conv_integer(x"40");
      PM_CAP_AUXCURRENT                                          : integer:= 0;
      PM_CAP_ID                                                  : integer:= conv_integer(x"01");
      PM_CAP_ON                                                  : string:= "TRUE";
      PM_CAP_PME_CLOCK                                           : string:= "FALSE";
      PM_CAP_RSVD_04                                             : integer:= 0;
      PM_CAP_VERSION                                             : integer:= 3;
      PM_CSR_BPCCEN                                              : string:= "FALSE";
      PM_CSR_B2B3                                                : string:= "FALSE";

      RECRC_CHK                                                  : integer:= 0;
      RECRC_CHK_TRIM                                             : string:= "FALSE";
      SELECT_DLL_IF                                              : string:= "FALSE";
      SPARE_BIT1                                                 : integer:= 0;
      SPARE_BIT2                                                 : integer:= 0;
      SPARE_BIT3                                                 : integer:= 0;
      SPARE_BIT4                                                 : integer:= 0;
      SPARE_BIT5                                                 : integer:= 0;
      SPARE_BIT6                                                 : integer:= 0;
      SPARE_BIT7                                                 : integer:= 0;
      SPARE_BIT8                                                 : integer:= 0;
      SPARE_BYTE0                                                : integer:= conv_integer(x"00");
      SPARE_BYTE1                                                : integer:= conv_integer(x"00");
      SPARE_BYTE2                                                : integer:= conv_integer(x"00");
      SPARE_BYTE3                                                : integer:= conv_integer(x"00");
      SPARE_WORD0                                                : integer:= conv_integer(x"00000000");
      SPARE_WORD1                                                : integer:= conv_integer(x"00000000");
      SPARE_WORD2                                                : integer:= conv_integer(x"00000000");
      SPARE_WORD3                                                : integer:= conv_integer(x"00000000");

      TL_RBYPASS                                                 : string:= "FALSE";
      TL_TFC_DISABLE                                             : string:= "FALSE";
      TL_TX_CHECKS_DISABLE                                       : string:= "FALSE";
      EXIT_LOOPBACK_ON_EI                                        : string:= "TRUE";
      UR_INV_REQ                                                 : string:= "TRUE";

      VC_CAP_ID                                                  : integer:= conv_integer(x"0002");
      VC_CAP_VERSION                                             : integer:= conv_integer(x"1");
      VSEC_CAP_HDR_ID                                            : integer:= conv_integer(x"1234");
      VSEC_CAP_HDR_LENGTH                                        : integer:= conv_integer(x"018");
      VSEC_CAP_HDR_REVISION                                      : integer:= conv_integer(x"1");
      VSEC_CAP_ID                                                : integer:= conv_integer(x"000b");
      VSEC_CAP_IS_LINK_VISIBLE                                   : string:= "TRUE";
      VSEC_CAP_VERSION                                           : integer:= conv_integer(x"1");

      C_BASEADDR_U                                               : integer:= conv_integer(x"FFFF");-- AXI Lite Base Address upper
      C_BASEADDR_L                                               : integer:= conv_integer(x"FFFF");-- AXI Lite Base Address lower
      C_HIGHADDR_U                                               : integer:= conv_integer(x"0000");-- AXI Lite High Address upper
      C_HIGHADDR_L                                               : integer:= conv_integer(x"0000");-- AXI Lite High Address lower
      C_MAX_LNK_WDT                                              : integer:= 1;                    -- Maximum Number of PCIE Lanes
      C_ROOT_PORT                                                : string:= "FALSE";               -- PCIe block is in root port mode
      C_RP_BAR_HIDE                                              : string:= "FALSE";               -- Hide RP PCIe BAR (prevent CPU from assigning address to RP BAR)
      C_RX_REALIGN                                               : string:= "TRUE";                -- Enable or Disable Realignment at RX Interface
      C_RX_PRESERVE_ORDER                                        : string:= "FALSE";               -- Preserve WR/ RD Ordering at the RX Interface
      C_LAST_CORE_CAP_ADDR                                       : integer:= conv_integer(x"000"); -- DWORD address of last enabled block capability
      C_VSEC_CAP_ADDR                                            : integer:= conv_integer(x"000"); -- DWORD address of start of VSEC Header
      C_VSEC_CAP_LAST                                            : string:= "FALSE";               -- VSEC next capability offset control
      C_VSEC_ID                                                  : integer:= conv_integer(x"0000");
      C_DEVICE_NUMBER                                            : integer:= 0;                    -- Device number for Root Port configurations only
      C_NUM_USER_INTR                                            : integer:= 0;                    -- Number of user interrupts in User interrupt vector
      C_USER_PTR                                                 : integer:= conv_integer(x"0000");-- Address pointer to User Space
      C_COMP_TIMEOUT                                             : integer:= 0;                    -- Completion Timout Value (0: 50us; 1:50ms)
      PTR_WIDTH                                                  : integer:= 4;
      C_FAMILY                                                   : string:= "V6";                  -- Targeted FPGA family

  --*******************************************************************
  -- S6 Parameter List
  --*******************************************************************

      USR_CFG                                                    : string:= "FALSE";
      USR_EXT_CFG                                                : string:= "FALSE";
      LINK_CAP_L0S_EXIT_LATENCY                                  : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY                                   : integer:= 7;
      PLM_AUTO_CONFIG                                            : string:= "FALSE";
      FAST_TRAIN                                                 : string:= "FALSE";
      PCIE_GENERIC                                               : integer:= conv_integer("000011101111");
      GTP_SEL                                                    : integer:= 0;
      CFG_VEN_ID                                                 : integer:= conv_integer(x"10EE");
      CFG_DEV_ID                                                 : integer:= conv_integer(x"0007");
      CFG_REV_ID                                                 : integer:= conv_integer(x"00");
      CFG_SUBSYS_VEN_ID                                          : integer:= conv_integer(x"10EE");
      CFG_SUBSYS_ID                                              : integer:= conv_integer(x"0007");

  --*******************************************************************
  -- K7 Parameter List
  --*******************************************************************

      AER_CAP_MULTIHEADER                                        : string:= "FALSE";
      AER_CAP_OPTIONAL_ERR_SUPPORT                               : integer:= conv_integer(x"000000");
      DEV_CAP2_ARI_FORWARDING_SUPPORTED                          : string:= "FALSE";
      DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED                    : string:= "FALSE";
      DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED                    : string:= "FALSE";
      DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED                        : string:= "FALSE";
      DEV_CAP2_CAS128_COMPLETER_SUPPORTED                        : string:= "FALSE";
      DEV_CAP2_TPH_COMPLETER_SUPPORTED                           : integer:= conv_integer(x"00");
      DEV_CONTROL_EXT_TAG_DEFAULT                                : string:= "FALSE";
      DISABLE_RX_POISONED_RESP                                   : string:= "FALSE";
      LINK_CAP_ASPM_OPTIONALITY                                  : string:= "FALSE";
      RBAR_BASE_PTR                                              : integer:= conv_integer(x"000");
      RBAR_CAP_CONTROL_ENCODEDBAR0                               : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR1                               : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR2                               : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR3                               : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR4                               : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR5                               : integer:= conv_integer(x"00");
      RBAR_CAP_INDEX0                                            : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX1                                            : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX2                                            : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX3                                            : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX4                                            : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX5                                            : integer:= conv_integer(x"0");
      RBAR_CAP_ON                                                : string:= "FALSE";
      RBAR_CAP_SUP0                                              : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP1                                              : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP2                                              : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP3                                              : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP4                                              : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP5                                              : integer:= conv_integer(x"00001");
      RBAR_NUM                                                   : integer:= conv_integer(x"0");
      TRN_NP_FC                                                  : string:= "TRUE";
      TRN_DW                                                     : string:= "FALSE";
      UR_ATOMIC                                                  : string:= "FALSE";
      UR_PRS_RESPONSE                                            : string:= "TRUE";
      USER_CLK2_DIV2                                             : string:= "FALSE";
      VC0_TOTAL_CREDITS_NPD                                      : integer:= 24;
      LINK_CAP_RSVD_23                                           : integer:= 0;
      CFG_ECRC_ERR_CPLSTAT                                       : integer:= 0;
      DISABLE_ERR_MSG                                            : string:= "FALSE";
      DISABLE_LOCKED_FILTER                                      : string:= "FALSE";
      DISABLE_PPM_FILTER                                         : string:= "FALSE";
      ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED                     : string:= "FALSE";
      INTERRUPT_STAT_AUTO                                        : string:= "TRUE";
      MPS_FORCE                                                  : string:= "FALSE";
      PM_ASPML0S_TIMEOUT                                         : integer:= conv_integer(x"0000");
      PM_ASPML0S_TIMEOUT_EN                                      : string:= "FALSE";
      PM_ASPML0S_TIMEOUT_FUNC                                    : integer:= 0;
      PM_ASPM_FASTEXIT                                           : string:= "FALSE";
      PM_MF                                                      : string:= "FALSE";
      RP_AUTO_SPD                                                : integer:= conv_integer(x"1");
      RP_AUTO_SPD_LOOPCNT                                        : integer:= conv_integer(x"1f");
      SIM_VERSION                                                : string:= "1.0";
      SSL_MESSAGE_AUTO                                           : string:= "FALSE";
      TECRC_EP_INV                                               : string:= "FALSE";
      UR_CFG1                                                    : string:= "TRUE";
      USE_RID_PINS                                               : string:= "FALSE";
      DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED                       : string:= "FALSE";
      DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED                      : string:= "FALSE";
      DEV_CAP2_LTR_MECHANISM_SUPPORTED                           : string:= "FALSE";
      DEV_CAP2_MAX_ENDEND_TLP_PREFIXES                           : integer:= conv_integer(x"0");
      DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING                        : string:= "FALSE";
      RBAR_CAP_ID                                                : integer:= conv_integer(x"0015");
      RBAR_CAP_NEXTPTR                                           : integer:= conv_integer(x"000");
      RBAR_CAP_VERSION                                           : integer:= conv_integer(x"1");
      PCIE_USE_MODE                                              : string:= "1.0";
      PCIE_GT_DEVICE                                             : string:= "GTP";
      PCIE_CHAN_BOND                                             : integer:= 1;
      PCIE_PLL_SEL                                               : string:= "CPLL";
      PCIE_ASYNC_EN                                              : string:= "FALSE";
      PCIE_TXBUF_EN                                              : string:= "FALSE";
      NO_SLV_ERR                    : string:= "FALSE";
      EXT_PIPE_INTERFACE                                         : string:= "FALSE"
   );
   port(
      -- 1. PCI Express (pci_exp) Interface
      ---------------------------------------------------------
      -- Tx
      pci_exp_txp                              : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      pci_exp_txn                              : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      -- Rx
      pci_exp_rxp                              : in  std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      pci_exp_rxn                              : in  std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);

qpll_drp_crscode	: in std_logic_vector(11 downto 0);
qpll_drp_fsm		: in std_logic_vector(17 downto 0);
qpll_drp_done     	: in std_logic_vector(1 downto 0);
qpll_drp_reset    	: in std_logic_vector(1 downto 0);       
qpll_qplllock    	: in std_logic_vector(1 downto 0);
qpll_qplloutclk    	: in std_logic_vector(1 downto 0);
qpll_qplloutrefclk	: in std_logic_vector(1 downto 0);
 qpll_qplld    : out std_logic_vector(1 downto 0)    ;
 qpll_qpllreset: out std_logic_vector(1 downto 0)    ;
 qpll_drp_clk: out std_logic_vector(1 downto 0)     ;
 qpll_drp_rst_n: out std_logic_vector(1 downto 0)     ;
 qpll_drp_ovrd: out std_logic_vector(1 downto 0)     ;
 qpll_drp_gen3: out std_logic_vector(1 downto 0)     ;
 qpll_drp_start: out std_logic_vector(1 downto 0)     ;

 pipe_txprbssel		:in std_logic_vector(2 downto 0);	
 pipe_rxprbssel	    	:in std_logic_vector(2 downto 0);    
 pipe_txprbsforceerr	:in std_logic;	
 pipe_rxprbscntreset	:in std_logic;	
 pipe_loopback 	    	:in std_logic_vector(2 downto 0);
 pipe_txinhibit               :in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);

 pipe_rxprbserr : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);


 pipe_rst_fsm 	:out std_logic_vector(4 downto 0);
 pipe_qrst_fsm	:out std_logic_vector(11 downto 0);	
 pipe_rate_fsm	:out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*5)-1 downto 0);	
 pipe_sync_fsm_tx	:out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*6)-1 downto 0);	
 pipe_sync_fsm_rx	:out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*7)-1 downto 0);	
 pipe_drp_fsm		:out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*7)-1 downto 0);	

 pipe_rst_idle	:out std_logic;	
 pipe_qrst_idle	:out std_logic;	
 pipe_rate_idle	:out std_logic;	
 pipe_eyescandataerror	:out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_rxstatus : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*3)-1 downto 0);    
 pipe_dmonitorout : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*15)-1 downto 0);

 pipe_cpll_lock          : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0); 
 pipe_qpll_lock          : out std_logic_vector(((LINK_CAP_MAX_LINK_WIDTH/8)+1)-1 downto 0); 
 pipe_rxpmaresetdone     : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);  
 pipe_rxbufstatus        : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*3)-1 downto 0);     
 pipe_txphaligndone      : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);   
 pipe_txphinitdone       : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);      
 pipe_txdlysresetdone    : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);    
 pipe_rxphaligndone      : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);     
 pipe_rxdlysresetdone    : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);      
 pipe_rxsyncdone         : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);      
 pipe_rxdisperr          : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*8)-1 downto 0);     
 pipe_rxnotintable       : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*8)-1 downto 0);     
 pipe_rxcommadet         : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);   

 gt_ch_drp_rdy	:out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	
 pipe_debug_0 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_1 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_2 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_3 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_4 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_5 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_6 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_7 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_8 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug_9 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 pipe_debug	:out std_logic_vector(31 downto 0);

 common_commands_in:in std_logic_vector(11 downto 0); 	
 pipe_rx_0_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_1_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_2_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_3_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_4_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_5_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_6_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_7_sigs	   :in std_logic_vector(24 downto 0);     
                          
 common_commands_out:out std_logic_vector(11 downto 0);	
 pipe_tx_0_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_1_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_2_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_3_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_4_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_5_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_6_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_7_sigs	    :out std_logic_vector(24 downto 0);    

 INT_PCLK_OUT_SLAVE	: out std_logic;	 
 INT_RXUSRCLK_OUT    	: out std_logic;   	
 INT_DCLK_OUT        	: out std_logic;   	
 INT_USERCLK1_OUT    	: out std_logic;   	
 INT_USERCLK2_OUT    	: out std_logic;   	
 INT_OOBCLK_OUT      	: out std_logic;   	
 INT_MMCM_LOCK_OUT   	: out std_logic;   	
 INT_QPLLLOCK_OUT	: out std_logic_vector(1 downto 0);	
 INT_QPLLOUTCLK_OUT	: out std_logic_vector(1 downto 0);	
 INT_QPLLOUTREFCLK_OUT	: out std_logic_vector(1 downto 0);	
 INT_RXOUTCLK_OUT 	: out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	      
 INT_PCLK_SEL_SLAVE	: in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	


    -------------Channel DRP---------------------------------
 ext_ch_gt_drpclk	 : out std_logic;	
 ext_ch_gt_drpaddr	 : in std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*9)-1 downto 0);	
 ext_ch_gt_drpen	 : in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	
 ext_ch_gt_drpdi	 : in std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*16)-1 downto 0);	
 ext_ch_gt_drpwe	 : in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	

 ext_ch_gt_drpdo	: out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*16)-1 downto 0);	
 ext_ch_gt_drprdy	: out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	
      ---------------------------------------------------------
      -- 2. Transaction (TRN) Interface
      ---------------------------------------------------------
      -- Rx
      rx_np_ok                                 : in  std_logic;
      rx_np_req                                : in  std_logic;

      ---------------------------------------------
      -- AXI TX - RW Interface
      -----------
      s_axis_rw_tdata                          : in  std_logic_vector(C_DATA_WIDTH-1 downto 0); -- RW data from user
      s_axis_rw_tvalid                         : in  std_logic;                                 -- RW data is valid
      s_axis_rw_tready                         : out std_logic;                                 -- RW ready for data
      s_axis_rw_tstrb                          : in  std_logic_vector(STRB_WIDTH-1 downto 0);   -- RW strobe byte enables
      s_axis_rw_tlast                          : in  std_logic;                                 -- RW data is last
      s_axis_rw_tuser                          : in  std_logic_vector(3 downto 0);              -- RW user signals

      -- AXI TX - RR Interface
      -------------
      s_axis_rr_tdata                          : in  std_logic_vector(C_DATA_WIDTH-1 downto 0); -- RR data from user
      s_axis_rr_tvalid                         : in  std_logic;                                 -- RR data is valid
      s_axis_rr_tready                         : out std_logic;                                 -- RR ready for data
      s_axis_rr_tstrb                          : in  std_logic_vector(STRB_WIDTH-1 downto 0);   -- RR strobe byte enables
      s_axis_rr_tlast                          : in  std_logic;                                 -- RR data is last
      s_axis_rr_tuser                          : in  std_logic_vector(3 downto 0);              -- RR user signals

      -- AXI TX - CC Interface
      -------------
      s_axis_cc_tdata                          : in  std_logic_vector(C_DATA_WIDTH-1 downto 0); -- CC data from user
      s_axis_cc_tvalid                         : in  std_logic;                                 -- CC data is valid
      s_axis_cc_tready                         : out std_logic;                                 -- CC ready for data
      s_axis_cc_tstrb                          : in  std_logic_vector(STRB_WIDTH-1 downto 0);   -- CC strobe byte enables
      s_axis_cc_tlast                          : in  std_logic;                                 -- CC data is last
      s_axis_cc_tuser                          : in  std_logic_vector(3 downto 0);              -- CC user signals

      -- AXI RX - CW Interface
      -------------
      m_axis_cw_tdata                          : out std_logic_vector(C_DATA_WIDTH-1 downto 0); -- CW data to user
      m_axis_cw_tvalid                         : out std_logic;                                 -- CW data is valid
      m_axis_cw_tready                         : in  std_logic;                                 -- CW ready for data
      m_axis_cw_tstrb                          : out std_logic_vector(STRB_WIDTH-1 downto 0);   -- CW strobe byte enables
      m_axis_cw_tlast                          : out std_logic;                                 -- CW data is last
      m_axis_cw_tuser                          : out std_logic_vector(21 downto 0);             -- CW user signals
 
      -- AXI RX - CR Interface
      -------------
      m_axis_cr_tdata                          : out std_logic_vector(C_DATA_WIDTH-1 downto 0); -- CR data to user
      m_axis_cr_tvalid                         : out std_logic;                                 -- CR data is valid
      m_axis_cr_tready                         : in  std_logic;                                 -- CR ready for data
      m_axis_cr_tstrb                          : out std_logic_vector(STRB_WIDTH-1 downto 0);   -- CR strobe byte enables
      m_axis_cr_tlast                          : out std_logic;                                 -- CR data is last
      m_axis_cr_tuser                          : out std_logic_vector(21 downto 0);             -- CR user signals

      -- AXI RX - RC Interface
      -------------
      m_axis_rc_tdata                          : out std_logic_vector(C_DATA_WIDTH-1 downto 0); -- RC data to user
      m_axis_rc_tvalid                         : out std_logic;                                 -- RC data is valid
      m_axis_rc_tready                         : in  std_logic;                                 -- RC ready for data
      m_axis_rc_tstrb                          : out std_logic_vector(STRB_WIDTH-1 downto 0);   -- RC strobe byte enables
      m_axis_rc_tlast                          : out std_logic;                                 -- RC data is last
      m_axis_rc_tuser                          : out std_logic_vector(21 downto 0);             -- RC user signals

      -- AXI -Lite Interface - CFG Block
      ---------------------------
      s_axi_ctl_awaddr                         : in  std_logic_vector(31 downto 0);             -- AXI Lite Write address
      s_axi_ctl_awvalid                        : in  std_logic;                                 -- AXI Lite Write Address Valid
      s_axi_ctl_awready                        : out std_logic;                                 -- AXI Lite Write Address Core ready
      s_axi_ctl_wdata                          : in  std_logic_vector(31 downto 0);             -- AXI Lite Write Data
      s_axi_ctl_wstrb                          : in  std_logic_vector(3 downto 0);              -- AXI Lite Write Data strobe
      s_axi_ctl_wvalid                         : in  std_logic;                                 -- AXI Lite Write data Valid
      s_axi_ctl_wready                         : out std_logic;                                 -- AXI Lite Write Data Core ready
      s_axi_ctl_bresp                          : out std_logic_vector(1 downto 0);              -- AXI Lite Write Data strobe
      s_axi_ctl_bvalid                         : out std_logic;                                 -- AXI Lite Write data Valid
      s_axi_ctl_bready                         : in  std_logic;                                 -- AXI Lite Write Data Core ready

      s_axi_ctl_araddr                         : in  std_logic_vector(31 downto 0);             -- AXI Lite Read address
      s_axi_ctl_arvalid                        : in  std_logic;                                 -- AXI Lite Read Address Valid
      s_axi_ctl_arready                        : out std_logic;                                 -- AXI Lite Read Address Core ready
      s_axi_ctl_rdata                          : out std_logic_vector(31 downto 0);             -- AXI Lite Read Data
      s_axi_ctl_rresp                          : out std_logic_vector(1 downto 0);              -- AXI Lite Read Data strobe
      s_axi_ctl_rvalid                         : out std_logic;                                 -- AXI Lite Read data Valid
      s_axi_ctl_rready                         : in  std_logic;                                 -- AXI Lite Read Data Core ready

      -- AXI Lite User IPIC Signals
      -----------------------------
      Bus2IP_CS                                : out std_logic;                                 -- Chip Select
      Bus2IP_BE                                : out std_logic_vector(3 downto 0);              -- Byte Enable Vector
      Bus2IP_RNW                               : out std_logic;                                 -- Read Npt Write Qualifier
      Bus2IP_Addr                              : out std_logic_vector(31 downto 0);             -- Address Bus
      Bus2IP_Data                              : out std_logic_vector(31 downto 0);             -- Write Data Bus
      IP2Bus_RdAck                             : in  std_logic;                                 -- Read Acknowledgement
      IP2Bus_WrAck                             : in  std_logic;                                 -- Write Acknowledgement
      IP2Bus_Data                              : in  std_logic_vector(31 downto 0);             -- Read Data Bus
      IP2Bus_Error                             : in  std_logic;                                 -- Error Qualifier

      --Interrupts
      -------------------
      ctl_intr                                 : out std_logic;                                 -- user interrupt
      ctl_user_intr                            : in  std_logic_vector(C_NUM_USER_INTR-1 downto 0);-- User interrupt vector used only in axi_pcie_mm_s
  
      -- User Misc.
      -------------
      --user_turnoff_ok                          : in  std_logic;                                 -- Turnoff OK from user
      --user_tcfg_gnt                            : in  std_logic;                                 -- Send cfg OK from user

      np_cpl_pending                           : in  std_logic;
      RP_bridge_en                             : out std_logic;

      ---------------------------------------------------------
      -- 3. Configuration (CFG) Interface
      ---------------------------------------------------------

      blk_err_cor                              : in  std_logic;
      blk_err_ur                               : in  std_logic;
      blk_err_ecrc                             : in  std_logic;
      blk_err_cpl_timeout                      : in  std_logic;
      blk_err_cpl_abort                        : in  std_logic;
      blk_err_cpl_unexpect                     : in  std_logic;
      blk_err_posted                           : in  std_logic;
      blk_err_locked                           : in  std_logic;
      blk_err_tlp_cpl_header                   : in  std_logic_vector(47 downto 0);
      blk_err_cpl_rdy                          : out std_logic;
      blk_interrupt                            : in  std_logic;
      blk_interrupt_rdy                        : out std_logic;
      blk_interrupt_assert                     : in  std_logic;
      blk_interrupt_di                         : in  std_logic_vector(7 downto 0);
      cfg_interrupt_do                         : out std_logic_vector(7 downto 0);
      blk_interrupt_mmenable                   : out std_logic_vector(2 downto 0);
      blk_interrupt_msienable                  : out std_logic;
      blk_interrupt_msixenable                 : out std_logic;
      blk_interrupt_msixfm                     : out std_logic;
      blk_trn_pending                          : in  std_logic;
      cfg_pm_send_pme_to                       : in  std_logic;
      blk_status                               : out std_logic_vector(15 downto 0);
      blk_command                              : out std_logic_vector(15 downto 0);
      blk_dstatus                              : out std_logic_vector(15 downto 0);
      blk_dcommand                             : out std_logic_vector(15 downto 0);
      blk_lstatus                              : out std_logic_vector(15 downto 0);
      blk_lcommand                             : out std_logic_vector(15 downto 0);
      blk_dcommand2                            : out std_logic_vector(15 downto 0);
      blk_pcie_link_state                      : out std_logic_vector(2 downto 0);
      blk_dsn                                  : in  std_logic_vector(63 downto 0);
      blk_pmcsr_pme_en                         : out std_logic;
      blk_pmcsr_pme_status                     : out std_logic;
      blk_pmcsr_powerstate                     : out std_logic_vector(1 downto 0);

      cfg_msg_received                         : out std_logic;
      blk_msg_data                             : out std_logic_vector(15 downto 0);
      blk_msg_received_err_cor                 : out std_logic;
      blk_msg_received_err_non_fatal           : out std_logic;
      blk_msg_received_err_fatal               : out std_logic;
      blk_msg_received_pme_to_ack              : out std_logic;
      blk_msg_received_assert_inta             : out std_logic;
      blk_msg_received_assert_intb             : out std_logic;
      blk_msg_received_assert_intc             : out std_logic;
      blk_msg_received_assert_intd             : out std_logic;
      blk_msg_received_deassert_inta           : out std_logic;
      blk_msg_received_deassert_intb           : out std_logic;
      blk_msg_received_deassert_intc           : out std_logic;
      blk_msg_received_deassert_intd           : out std_logic;

      blk_link_up                              : out std_logic;

      blk_ds_bus_number                        : in  std_logic_vector(7 downto 0);
      blk_ds_device_number                     : in  std_logic_vector(4 downto 0);

      -- Only for End point Cores
      blk_to_turnoff                           : out  std_logic;
      blk_turnoff_ok                           : in std_logic;
      blk_pm_wake                              : in std_logic;

      blk_bus_number                           : out std_logic_vector(7 downto 0);
      blk_device_number                        : out std_logic_vector(4 downto 0);
      blk_function_number                      : out std_logic_vector(2 downto 0);

      ---------------------------------------------------------
      -- 4. Physical Layer Control and Status (PL) Interface
      ---------------------------------------------------------

      blk_pl_initial_link_width                : out std_logic_vector(2 downto 0);
      blk_pl_lane_reversal_mode                : out std_logic_vector(1 downto 0);
      blk_pl_link_gen2_capable                 : out std_logic;
      blk_pl_link_partner_gen2_supported       : out std_logic;
      blk_pl_link_upcfg_capable                : out std_logic;
      blk_pl_ltssm_state                       : out std_logic_vector(5 downto 0);
      blk_pl_sel_link_rate                     : out std_logic;
      blk_pl_sel_link_width                    : out std_logic_vector(1 downto 0);
      blk_pl_upstream_prefer_deemph            : in  std_logic;
      blk_pl_hot_rst                           : out std_logic;

      -- Flow Control
      blk_fc_cpld                              : out std_logic_vector(11 downto 0);
      blk_fc_cplh                              : out std_logic_vector(7 downto 0);
      blk_fc_npd                               : out std_logic_vector(11 downto 0);
      blk_fc_nph                               : out std_logic_vector(7 downto 0);
      blk_fc_pd                                : out std_logic_vector(11 downto 0);
      blk_fc_ph                                : out std_logic_vector(7 downto 0);
      blk_fc_sel                               : in  std_logic_vector(2 downto 0);

      -- Tx

      blk_tbuf_av                              : out std_logic_vector(5 downto 0);
      blk_tcfg_req                             : out std_logic;                                    
      blk_tcfg_gnt                             : in  std_logic;                               

      tx_err_drop                              : out std_logic;                     

      --S-6 Specific

      cfg_do                                   : out std_logic_vector(31 downto 0);
      cfg_rd_wr_done                           : out std_logic;                                
      cfg_dwaddr                               : in  std_logic_vector(9 downto 0);
      cfg_rd_en                                : in  std_logic;                          

      ---------------------------------------------------------
      -- 5. System  (SYS) Interface
      ---------------------------------------------------------

      com_sysclk                               : in  std_logic;
      com_sysrst                               : in  std_logic;
      mmcm_lock                                : out std_logic;
      com_iclk                                 : out std_logic;
      com_cclk                                 : out std_logic;
      com_corereset                            : out std_logic;

      clk_fab_refclk                           : in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      clk_pclk                                 : in std_logic;
      clk_rxusrclk                             : in std_logic;
      clk_dclk                                 : in std_logic;
      clk_userclk1                             : in std_logic;
      clk_userclk2                             : in std_logic;
      clk_oobclk_in                            : in std_logic;
      clk_mmcm_lock                            : in std_logic;
      clk_txoutclk                             : out std_logic;
      clk_rxoutclk                             : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      clk_pclk_sel                             : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      clk_gen3                                 : out std_logic;
      PIPE_MMCM_RST_N                          : in std_logic;
      config_gen_req                           : out std_logic
      
   );

end axi_enhanced_pcie;

architecture structure of axi_enhanced_pcie is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

component axi_pcie_v2_9_14_enhanced_core_top_wrap
   generic(
      C_DATA_WIDTH                             : integer:= 64;
      STRB_WIDTH                               : integer:= 8;
      BAR0_U                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR0_L                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR1_U                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR1_L                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR2_U                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR2_L                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR3_U                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR3_L                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR4_U                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR4_L                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR5_U                                   : std_logic_vector(15 downto 0):= x"ffff";
      BAR5_L                                   : std_logic_vector(15 downto 0):= x"ffff";

      CARDBUS_CIS_POINTER                      : integer:= conv_integer(x"00000000");
      CLASS_CODE                               : integer:= conv_integer(x"060000");
      CMD_INTX_IMPLEMENTED                     : string:= "TRUE";
      CPL_TIMEOUT_DISABLE_SUPPORTED            : string:= "FALSE";
      CPL_TIMEOUT_RANGES_SUPPORTED             : integer:= conv_integer(x"2");

      DEV_CAP_EXT_TAG_SUPPORTED                : string:= "FALSE";
      DEV_CAP_MAX_PAYLOAD_SUPPORTED            : integer:= 2;
      DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT        : integer:= 0;
      DEVICE_ID                                : integer:= conv_integer(x"6011");

      DISABLE_LANE_REVERSAL                    : string:= "TRUE";
      DISABLE_SCRAMBLING                       : string:= "FALSE";
      DSN_BASE_PTR                             : integer:= conv_integer(x"100");
      DSN_CAP_NEXTPTR                          : integer:= conv_integer(x"000");
      DSN_CAP_ON                               : string:= "TRUE";

      ENABLE_MSG_ROUTE                         : integer:= conv_integer(x"000");
      ENABLE_RX_TD_ECRC_TRIM                   : string:= "FALSE";
      EXPANSION_ROM_U                          : integer:= conv_integer(x"ffff");
      EXPANSION_ROM_L                          : integer:= conv_integer(x"f001");
      EXT_CFG_CAP_PTR                          : integer:= conv_integer(x"3f");
      EXT_CFG_XP_CAP_PTR                       : integer:= conv_integer(x"3ff");
      HEADER_TYPE                              : integer:= conv_integer(x"00");
      INTERRUPT_PIN                            : integer:= conv_integer(x"01");

      LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP   : string:= "FALSE";
      LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP : string:= "FALSE";
      LINK_CAP_MAX_LINK_SPEED                  : integer:= conv_integer(x"1");
      LINK_CAP_MAX_LINK_WIDTH                  : integer:= conv_integer(x"01");
      LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE     : string:= "FALSE";

      LINK_CONTROL_RCB                         : integer:= 0;
      LINK_CTRL2_DEEMPHASIS                    : string:= "FALSE";
      LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE   : string:= "FALSE";
      LINK_CTRL2_TARGET_LINK_SPEED             : integer:= conv_integer(x"0");
      LINK_STATUS_SLOT_CLOCK_CONFIG            : string:= "FALSE";

      LL_ACK_TIMEOUT                           : integer:= conv_integer(x"0000");
      LL_ACK_TIMEOUT_EN                        : string:= "FALSE";
      LL_ACK_TIMEOUT_FUNC                      : integer:= 0;
      LL_REPLAY_TIMEOUT                        : integer:= conv_integer(x"0026");
      LL_REPLAY_TIMEOUT_EN                     : string:= "TRUE";
      LL_REPLAY_TIMEOUT_FUNC                   : integer:= 1;

      LTSSM_MAX_LINK_WIDTH                     : integer:= conv_integer(x"1");
      MSI_DECODE_ENABLE                        : string:= "TRUE";
      MSI_CAP_MULTIMSGCAP                      : integer:= 0;
      MSI_CAP_MULTIMSG_EXTENSION               : integer:= 0;
      MSI_CAP_ON                               : string:= "TRUE";
      MSI_CAP_PER_VECTOR_MASKING_CAPABLE       : string:= "FALSE";
      MSI_CAP_64_BIT_ADDR_CAPABLE              : string:= "TRUE";

      MSIX_CAP_ON                              : string:= "FALSE";
      MSIX_CAP_PBA_BIR                         : integer:= 0;
      MSIX_CAP_PBA_OFFSET                      : integer:= conv_integer(x"00000000");
      MSIX_CAP_TABLE_BIR                       : integer:= 0;
      MSIX_CAP_TABLE_OFFSET                    : integer:= conv_integer(x"00000000");
      MSIX_CAP_TABLE_SIZE                      : integer:= conv_integer(x"000");

      PCIE_CAP_DEVICE_PORT_TYPE                : integer:= conv_integer(x"0");
      PCIE_CAP_INT_MSG_NUM                     : integer:= conv_integer(x"01");
      PCIE_CAP_NEXTPTR                         : integer:= conv_integer(x"00");
      PCIE_DRP_ENABLE                          : string:= "FALSE";
      PIPE_PIPELINE_STAGES                     : integer:= 0;  -- 0 - 0 stages, 1 - 1 stage, 2 - 2 stages

      PM_CAP_DSI                               : string:= "FALSE";
      PM_CAP_D1SUPPORT                         : string:= "FALSE";
      PM_CAP_D2SUPPORT                         : string:= "FALSE";
      PM_CAP_NEXTPTR                           : integer:= conv_integer(x"48");
      PM_CAP_PMESUPPORT                        : integer:= conv_integer(x"0f");
      PM_CSR_NOSOFTRST                         : string:= "TRUE";

      PM_DATA_SCALE0                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE1                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE2                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE3                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE4                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE5                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE6                           : integer:= conv_integer(x"0");
      PM_DATA_SCALE7                           : integer:= conv_integer(x"0");

      PM_DATA0                                 : integer:= conv_integer(x"00");
      PM_DATA1                                 : integer:= conv_integer(x"00");
      PM_DATA2                                 : integer:= conv_integer(x"00");
      PM_DATA3                                 : integer:= conv_integer(x"00");
      PM_DATA4                                 : integer:= conv_integer(x"00");
      PM_DATA5                                 : integer:= conv_integer(x"00");
      PM_DATA6                                 : integer:= conv_integer(x"00");
      PM_DATA7                                 : integer:= conv_integer(x"00");

      REF_CLK_FREQ                             : integer:= 0;  -- 0 - 100 MHz, 1 - 125 MHz, 2 - 250 MHz
      REVISION_ID                              : integer:= conv_integer(x"00");
      ROOT_CAP_CRS_SW_VISIBILITY               : string:= "FALSE";
      SPARE_BIT0                               : integer:= 0;
      SUBSYSTEM_ID                             : integer:= conv_integer(x"0007");
      SUBSYSTEM_VENDOR_ID                      : integer:= conv_integer(x"10ee");

      SLOT_CAP_ATT_BUTTON_PRESENT              : string:= "FALSE";
      SLOT_CAP_ATT_INDICATOR_PRESENT           : string:= "FALSE";
      SLOT_CAP_ELEC_INTERLOCK_PRESENT          : string:= "FALSE";
      SLOT_CAP_HOTPLUG_CAPABLE                 : string:= "FALSE";
      SLOT_CAP_HOTPLUG_SURPRISE                : string:= "FALSE";
      SLOT_CAP_MRL_SENSOR_PRESENT              : string:= "FALSE";
      SLOT_CAP_NO_CMD_COMPLETED_SUPPORT        : string:= "FALSE";
      SLOT_CAP_PHYSICAL_SLOT_NUM               : integer:= conv_integer(x"0000");
      SLOT_CAP_POWER_CONTROLLER_PRESENT        : string:= "FALSE";
      SLOT_CAP_POWER_INDICATOR_PRESENT         : string:= "FALSE";
      SLOT_CAP_SLOT_POWER_LIMIT_SCALE          : integer:= 0;
      SLOT_CAP_SLOT_POWER_LIMIT_VALUE          : integer:= conv_integer(x"00");

      TL_RX_RAM_RADDR_LATENCY                  : integer:= 0;
      TL_RX_RAM_RDATA_LATENCY                  : integer:= 2;
      TL_RX_RAM_WRITE_LATENCY                  : integer:= 0;
      TL_TX_RAM_RADDR_LATENCY                  : integer:= 0;
      TL_TX_RAM_RDATA_LATENCY                  : integer:= 2;
      TL_TX_RAM_WRITE_LATENCY                  : integer:= 0;

      UPCONFIG_CAPABLE                         : string:= "TRUE";
      UPSTREAM_FACING                          : STRING:= "FALSE";
      USER_CLK_FREQ                            : integer:= 1;--3
      VC_BASE_PTR                              : integer:= conv_integer(x"000");
      VC_CAP_NEXTPTR                           : integer:= conv_integer(x"000");
      VC_CAP_ON                                : string:= "FALSE";
      VC_CAP_REJECT_SNOOP_TRANSACTIONS         : string:= "FALSE";

      VC0_CPL_INFINITE                         : string:= "TRUE";
      VC0_RX_RAM_LIMIT                         : integer:= conv_integer(x"07ff");
      VC0_TOTAL_CREDITS_CD                     : integer:= 308;
      VC0_TOTAL_CREDITS_CH                     : integer:= 36;
      VC0_TOTAL_CREDITS_NPH                    : integer:= 12;
      VC0_TOTAL_CREDITS_PD                     : integer:= 308;
      VC0_TOTAL_CREDITS_PH                     : integer:= 32;
      VC0_TX_LASTPACKET                        : integer:= 29;

      VENDOR_ID                                : integer:= conv_integer(x"10ee");
      VSEC_BASE_PTR                            : integer:= conv_integer(x"000");
      VSEC_CAP_NEXTPTR                         : integer:= conv_integer(x"000");
      VSEC_CAP_ON                              : string:= "FALSE";

      ALLOW_X8_GEN2                            : string:= "FALSE";
      AER_BASE_PTR                             : integer:= conv_integer(x"128");
      AER_CAP_ECRC_CHECK_CAPABLE               : string:= "FALSE";
      AER_CAP_ECRC_GEN_CAPABLE                 : string:= "FALSE";
      AER_CAP_ID                               : integer:= conv_integer(x"0001");
      AER_CAP_INT_MSG_NUM_MSI                  : integer:= conv_integer(x"0a");
      AER_CAP_INT_MSG_NUM_MSIX                 : integer:= conv_integer(x"15");
      AER_CAP_NEXTPTR                          : integer:= conv_integer(x"160");
      AER_CAP_ON                               : string:= "FALSE";
      AER_CAP_PERMIT_ROOTERR_UPDATE            : string:= "TRUE";
      AER_CAP_VERSION                          : integer:= conv_integer(x"1");

      CAPABILITIES_PTR                         : integer:= conv_integer(x"40");
      CRM_MODULE_RSTS                          : integer:= conv_integer(x"00");
      DEV_CAP_ENDPOINT_L0S_LATENCY             : integer:= 0;
      DEV_CAP_ENDPOINT_L1_LATENCY              : integer:= 0;
      DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE     : string:= "FALSE";
      DEV_CAP_ROLE_BASED_ERROR                 : string:= "TRUE";
      DEV_CAP_RSVD_14_12                       : integer:= 0;
      DEV_CAP_RSVD_17_16                       : integer:= 0;
      DEV_CAP_RSVD_31_29                       : integer:= 0;
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE      : string:= "TRUE";
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE      : string:= "TRUE";
      DEV_CONTROL_AUX_POWER_SUPPORTED          : string:= "FALSE";

      DISABLE_ASPM_L1_TIMER                    : string:= "FALSE";
      DISABLE_BAR_FILTERING                    : string:= "FALSE";
      DISABLE_ID_CHECK                         : string:= "FALSE";
      DISABLE_RX_TC_FILTER                     : string:= "FALSE";
      DNSTREAM_LINK_NUM                        : integer:= conv_integer(x"00");

      DS_PORT_HOT_RST                          : string:= "FALSE";  -- FALSE - for ROOT PORT(default), TRUE - for DOWNSTREAM PORT 
      DSN_CAP_ID                               : integer:= conv_integer(x"0003");
      DSN_CAP_VERSION                          : integer:= conv_integer(x"1");
      ENTER_RVRY_EI_L0                         : string:= "TRUE";
      INFER_EI                                 : integer:= conv_integer(x"0c");
      IS_SWITCH                                : string:= "FALSE";

      LAST_CONFIG_DWORD                        : integer:= conv_integer(x"3ff");
      LINK_CAP_ASPM_SUPPORT                    : integer:= 1;
      LINK_CAP_CLOCK_POWER_MANAGEMENT          : string:= "FALSE";
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    : integer:= 7;
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    : integer:= 7;
      LINK_CAP_L0S_EXIT_LATENCY_GEN1           : integer:= 7;
      LINK_CAP_L0S_EXIT_LATENCY_GEN2           : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1     : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2     : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_GEN1            : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY_GEN2            : integer:= 7;
      LINK_CAP_RSVD_23_22                      : integer:= 0;

      MSI_BASE_PTR                             : integer:= conv_integer(x"48");
      MSI_CAP_ID                               : integer:= conv_integer(x"05");
      MSI_CAP_NEXTPTR                          : integer:= conv_integer(x"60");
      MSIX_BASE_PTR                            : integer:= conv_integer(x"9c");
      MSIX_CAP_ID                              : integer:= conv_integer(x"11");
      MSIX_CAP_NEXTPTR                         : integer:= conv_integer(x"00");
      N_FTS_COMCLK_GEN1                        : integer:= 255;
      N_FTS_COMCLK_GEN2                        : integer:= 254;
      N_FTS_GEN1                               : integer:= 255;
      N_FTS_GEN2                               : integer:= 255;

      PCIE_BASE_PTR                            : integer:= conv_integer(x"60");
      PCIE_CAP_CAPABILITY_ID                   : integer:= conv_integer(x"10");
      PCIE_CAP_CAPABILITY_VERSION              : integer:= conv_integer(x"2");
      PCIE_CAP_ON                              : string:= "TRUE";
      PCIE_CAP_RSVD_15_14                      : integer:= 0;
      PCIE_CAP_SLOT_IMPLEMENTED                : string:= "FALSE";
      PCIE_REVISION                            : integer:= 2;
      PGL0_LANE                                : integer:= 0;
      PGL1_LANE                                : integer:= 1;
      PGL2_LANE                                : integer:= 2;
      PGL3_LANE                                : integer:= 3;
      PGL4_LANE                                : integer:= 4;
      PGL5_LANE                                : integer:= 5;
      PGL6_LANE                                : integer:= 6;
      PGL7_LANE                                : integer:= 7;
      PL_AUTO_CONFIG                           : integer:= 0;
      PL_FAST_TRAIN                            : string:= "FALSE";
      PCIE_EXT_CLK                             : string:= "TRUE";
      NO_SLV_ERR                    : string:= "FALSE";
       PCIE_EXT_GT_COMMON : string:= "FALSE";
       EXT_CH_GT_DRP : string:= "FALSE";

 TX_MARGIN_FULL_0  :integer:= conv_integer (x"4F");
 TX_MARGIN_FULL_1  :integer:= conv_integer (x"4e");
 TX_MARGIN_FULL_2  :integer:= conv_integer (x"4d");
 TX_MARGIN_FULL_3  :integer:= conv_integer (x"4c");
 TX_MARGIN_FULL_4  :integer:= conv_integer (x"43");
 TX_MARGIN_LOW_0   :integer:= conv_integer (x"45");
 TX_MARGIN_LOW_1   :integer:= conv_integer (x"46");
 TX_MARGIN_LOW_2   :integer:= conv_integer (x"43");
 TX_MARGIN_LOW_3   :integer:= conv_integer (x"42");
 TX_MARGIN_LOW_4   :integer:=conv_integer  (x"40");
      PM_BASE_PTR                              : integer:= conv_integer(x"40");
      PM_CAP_AUXCURRENT                        : integer:= 0;
      PM_CAP_ID                                : integer:= conv_integer(x"01");
      PM_CAP_ON                                : string:= "TRUE";
      PM_CAP_PME_CLOCK                         : string:= "FALSE";
      PM_CAP_RSVD_04                           : integer:= 0;
      PM_CAP_VERSION                           : integer:= 3;
      PM_CSR_BPCCEN                            : string:= "FALSE";
      PM_CSR_B2B3                              : string:= "FALSE";

      RECRC_CHK                                : integer:= 0;
      RECRC_CHK_TRIM                           : string:= "FALSE";
      SELECT_DLL_IF                            : string:= "FALSE";
      SPARE_BIT1                               : integer:= 0;
      SPARE_BIT2                               : integer:= 0;
      SPARE_BIT3                               : integer:= 0;
      SPARE_BIT4                               : integer:= 0;
      SPARE_BIT5                               : integer:= 0;
      SPARE_BIT6                               : integer:= 0;
      SPARE_BIT7                               : integer:= 0;
      SPARE_BIT8                               : integer:= 0;
      SPARE_BYTE0                              : integer:= conv_integer(x"00");
      SPARE_BYTE1                              : integer:= conv_integer(x"00");
      SPARE_BYTE2                              : integer:= conv_integer(x"00");
      SPARE_BYTE3                              : integer:= conv_integer(x"00");
      SPARE_WORD0                              : integer:= conv_integer(x"00000000");
      SPARE_WORD1                              : integer:= conv_integer(x"00000000");
      SPARE_WORD2                              : integer:= conv_integer(x"00000000");
      SPARE_WORD3                              : integer:= conv_integer(x"00000000");

      TL_RBYPASS                               : string:= "FALSE";
      TL_TFC_DISABLE                           : string:= "FALSE";
      TL_TX_CHECKS_DISABLE                     : string:= "FALSE";
      EXIT_LOOPBACK_ON_EI                      : string:= "TRUE";
      UR_INV_REQ                               : string:= "TRUE";

      VC_CAP_ID                                : integer:= conv_integer(x"0002");
      VC_CAP_VERSION                           : integer:= conv_integer(x"1");
      VSEC_CAP_HDR_ID                          : integer:= conv_integer(x"1234");
      VSEC_CAP_HDR_LENGTH                      : integer:= conv_integer(x"018");
      VSEC_CAP_HDR_REVISION                    : integer:= conv_integer(x"1");
      VSEC_CAP_ID                              : integer:= conv_integer(x"000b");
      VSEC_CAP_IS_LINK_VISIBLE                 : string:= "TRUE";
      VSEC_CAP_VERSION                         : integer:= conv_integer(x"1");

      C_BASEADDR_U                             : integer:= conv_integer(x"FFFF");-- AXI Lite Base Address upper
      C_BASEADDR_L                             : integer:= conv_integer(x"FFFF");-- AXI Lite Base Address lower
      C_HIGHADDR_U                             : integer:= conv_integer(x"0000");-- AXI Lite High Address upper
      C_HIGHADDR_L                             : integer:= conv_integer(x"0000");-- AXI Lite High Address lower

      C_MAX_LNK_WDT                            : integer:= 1;                    -- Maximum Number of PCIE Lanes
      C_ROOT_PORT                              : string:= "FALSE";               -- PCIe block is in root port mode
      C_RP_BAR_HIDE                            : string:= "FALSE";               -- Hide RP PCIe BAR (prevent CPU from assigning address to RP BAR)
      C_RX_REALIGN                             : string:= "TRUE";                -- Enable or Disable Realignment at RX Interface
      C_RX_PRESERVE_ORDER                      : string:= "FALSE";               -- Preserve WR/ RD Ordering at the RX Interface
      C_LAST_CORE_CAP_ADDR                     : integer:= conv_integer(x"000"); -- DWORD address of last enabled block capability
      C_VSEC_CAP_ADDR                          : integer:= conv_integer(x"000"); -- DWORD address of start of VSEC Header
      C_VSEC_CAP_LAST                          : string:= "FALSE";               -- VSEC next capability offset control
      C_VSEC_ID                                : integer:= conv_integer(x"0000");
      C_DEVICE_NUMBER                          : integer:= 0;                    -- Device number for Root Port configurations only
      C_NUM_USER_INTR                          : integer:= 0;                    -- Number of user interrupts in User interrupt vector
      C_USER_PTR                               : integer:= conv_integer(x"0000"); -- Address pointer to User Space
      C_COMP_TIMEOUT                           : integer:= 0;                    -- Completion Timout Value (0: 50us; 1:50ms)
      PTR_WIDTH                                : integer:= 4;
      C_FAMILY                                 : string:= "V6";                   -- Targeted FPGA family

  --*******************************************************************
  -- S6 Parameter List
  --*******************************************************************

      USR_CFG                                  : string:= "FALSE";
      USR_EXT_CFG                              : string:= "FALSE";
      LINK_CAP_L0S_EXIT_LATENCY                : integer:= 7;
      LINK_CAP_L1_EXIT_LATENCY                 : integer:= 7;
      PLM_AUTO_CONFIG                          : string:= "FALSE";
      FAST_TRAIN                               : string:= "FALSE";
      PCIE_GENERIC                             : integer:= conv_integer("000011101111");
      GTP_SEL                                  : integer:= 0;
      CFG_VEN_ID                               : integer:= conv_integer(x"10EE");
      CFG_DEV_ID                               : integer:= conv_integer(x"0007");
      CFG_REV_ID                               : integer:= conv_integer(x"00");
      CFG_SUBSYS_VEN_ID                        : integer:= conv_integer(x"10EE");
      CFG_SUBSYS_ID                            : integer:= conv_integer(x"0007");

  --*******************************************************************
  -- K7 Parameter List
  --*******************************************************************

      AER_CAP_MULTIHEADER                      : string:= "FALSE";
      AER_CAP_OPTIONAL_ERR_SUPPORT             : integer:= conv_integer(x"000000");
      DEV_CAP2_ARI_FORWARDING_SUPPORTED        : string:= "FALSE";
      DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED  : string:= "FALSE";
      DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED  : string:= "FALSE";
      DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED      : string:= "FALSE";
      DEV_CAP2_CAS128_COMPLETER_SUPPORTED      : string:= "FALSE";
      DEV_CAP2_TPH_COMPLETER_SUPPORTED         : integer:= conv_integer(x"00");
      DEV_CONTROL_EXT_TAG_DEFAULT              : string:= "FALSE";
      DISABLE_RX_POISONED_RESP                 : string:= "FALSE";
      LINK_CAP_ASPM_OPTIONALITY                : string:= "FALSE";
      RBAR_BASE_PTR                            : integer:= conv_integer(x"000");
      RBAR_CAP_CONTROL_ENCODEDBAR0             : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR1             : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR2             : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR3             : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR4             : integer:= conv_integer(x"00");
      RBAR_CAP_CONTROL_ENCODEDBAR5             : integer:= conv_integer(x"00");
      RBAR_CAP_INDEX0                          : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX1                          : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX2                          : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX3                          : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX4                          : integer:= conv_integer(x"0");
      RBAR_CAP_INDEX5                          : integer:= conv_integer(x"0");
      RBAR_CAP_ON                              : string:= "FALSE";
      RBAR_CAP_SUP0                            : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP1                            : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP2                            : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP3                            : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP4                            : integer:= conv_integer(x"00001");
      RBAR_CAP_SUP5                            : integer:= conv_integer(x"00001");
      RBAR_NUM                                 : integer:= conv_integer(x"0");
      TRN_NP_FC                                : string:= "TRUE";
      TRN_DW                                   : string:= "FALSE";
      UR_ATOMIC                                : string:= "FALSE";
      UR_PRS_RESPONSE                          : string:= "TRUE";
      USER_CLK2_DIV2                           : string:= "FALSE";
      VC0_TOTAL_CREDITS_NPD                    : integer:= 24;
      LINK_CAP_RSVD_23                         : integer:= 0;
      CFG_ECRC_ERR_CPLSTAT                     : integer:= 0;
      DISABLE_ERR_MSG                          : string:= "FALSE";
      DISABLE_LOCKED_FILTER                    : string:= "FALSE";
      DISABLE_PPM_FILTER                       : string:= "FALSE";
      ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED   : string:= "FALSE";
      INTERRUPT_STAT_AUTO                      : string:= "TRUE";
      MPS_FORCE                                : string:= "FALSE";
      PM_ASPML0S_TIMEOUT                       : integer:= conv_integer(x"0000");
      PM_ASPML0S_TIMEOUT_EN                    : string:= "FALSE";
      PM_ASPML0S_TIMEOUT_FUNC                  : integer:= 0;
      PM_ASPM_FASTEXIT                         : string:= "FALSE";
      PM_MF                                    : string:= "FALSE";
      RP_AUTO_SPD                              : integer:= conv_integer(x"1");
      RP_AUTO_SPD_LOOPCNT                      : integer:= conv_integer(x"1f");
      SIM_VERSION                              : string:= "1.0";
      SSL_MESSAGE_AUTO                         : string:= "FALSE";
      TECRC_EP_INV                             : string:= "FALSE";
      UR_CFG1                                  : string:= "TRUE";
      USE_RID_PINS                             : string:= "FALSE";
      DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED     : string:= "FALSE";
      DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED    : string:= "FALSE";
      DEV_CAP2_LTR_MECHANISM_SUPPORTED         : string:= "FALSE";
      DEV_CAP2_MAX_ENDEND_TLP_PREFIXES         : integer:= conv_integer(x"0");
      DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING      : string:= "FALSE";
      RBAR_CAP_ID                              : integer:= conv_integer(x"0015");
      RBAR_CAP_NEXTPTR                         : integer:= conv_integer(x"000");
      RBAR_CAP_VERSION                         : integer:= conv_integer(x"1");
      PCIE_USE_MODE                            : string:= "1.0";
      PCIE_GT_DEVICE                           : string:= "GTP";
      PCIE_CHAN_BOND                           : integer:= 1;
      PCIE_PLL_SEL                             : string:= "CPLL";
      PCIE_ASYNC_EN                            : string:= "FALSE";
      PCIE_TXBUF_EN                            : string:= "FALSE";
      EXT_PIPE_INTERFACE                       : string:= "FALSE"
   );
   port(
      -- 1. PCI Express (pci_exp) Interface
      ---------------------------------------------------------
      -- Tx
      pci_exp_txp                              : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      pci_exp_txn                              : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      -- Rx
      pci_exp_rxp                              : in  std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      pci_exp_rxn                              : in  std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
 qpll_drp_crscode      : in std_logic_vector(11 downto 0);
 qpll_drp_fsm          : in std_logic_vector(17 downto 0);
 qpll_drp_done         : in std_logic_vector(1 downto 0);
 qpll_drp_reset        : in std_logic_vector(1 downto 0);
 qpll_qplllock         : in std_logic_vector(1 downto 0);
 qpll_qplloutclk       : in std_logic_vector(1 downto 0);
 qpll_qplloutrefclk    : in std_logic_vector(1 downto 0);
 qpll_qplld    : out std_logic_vector(1 downto 0)    ;
  qpll_qpllreset: out std_logic_vector(1 downto 0)    ;
  qpll_drp_clk: out std_logic_vector(1 downto 0)     ;
  qpll_drp_rst_n: out std_logic_vector(1 downto 0)     ;
  qpll_drp_ovrd: out std_logic_vector(1 downto 0)     ;
  qpll_drp_gen3: out std_logic_vector(1 downto 0)     ;
  qpll_drp_start: out std_logic_vector(1 downto 0)     ;

  pipe_txprbssel               :in std_logic_vector(2 downto 0);
  pipe_rxprbssel               :in std_logic_vector(2 downto 0);
  pipe_txprbsforceerr  :in std_logic;
  pipe_rxprbscntreset  :in std_logic;
  pipe_loopback                :in std_logic_vector(2 downto 0);
  pipe_txinhibit               :in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);

  pipe_rxprbserr : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);


  pipe_rst_fsm         :out std_logic_vector(4 downto 0);
  pipe_qrst_fsm        :out std_logic_vector(11 downto 0);
  pipe_rate_fsm        :out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*5)-1 downto 0);
  pipe_sync_fsm_tx     :out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*6)-1 downto 0);
  pipe_sync_fsm_rx     :out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*7)-1 downto 0);
  pipe_drp_fsm         :out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*7)-1 downto 0);

  pipe_rst_idle        :out std_logic;
  pipe_qrst_idle       :out std_logic;
  pipe_rate_idle       :out std_logic;
  pipe_eyescandataerror	:out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_rxstatus : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*3)-1 downto 0);    
  pipe_dmonitorout : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*15)-1 downto 0);

  pipe_cpll_lock          : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0); 
  pipe_qpll_lock          : out std_logic_vector(((LINK_CAP_MAX_LINK_WIDTH/8)+1)-1 downto 0); 
  pipe_rxpmaresetdone     : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);  
  pipe_rxbufstatus        : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*3)-1 downto 0);     
  pipe_txphaligndone      : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);   
  pipe_txphinitdone       : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);      
  pipe_txdlysresetdone    : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);    
  pipe_rxphaligndone      : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);     
  pipe_rxdlysresetdone    : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);      
  pipe_rxsyncdone         : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);      
  pipe_rxdisperr          : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*8)-1 downto 0);     
  pipe_rxnotintable       : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*8)-1 downto 0);     
  pipe_rxcommadet         : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);   

  gt_ch_drp_rdy        :out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_0 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_1 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_2 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_3 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_4 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_5 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_6 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_7 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_8 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug_9 : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  pipe_debug   :out std_logic_vector(31 downto 0);

 common_commands_in:in std_logic_vector(11 downto 0); 	
 pipe_rx_0_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_1_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_2_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_3_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_4_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_5_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_6_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_7_sigs	   :in std_logic_vector(24 downto 0);     
                          
 common_commands_out:out std_logic_vector(11 downto 0);	
 pipe_tx_0_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_1_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_2_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_3_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_4_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_5_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_6_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_7_sigs	    :out std_logic_vector(24 downto 0);    

 INT_PCLK_OUT_SLAVE	: out std_logic;	 
 INT_RXUSRCLK_OUT    	: out std_logic;   	
 INT_DCLK_OUT        	: out std_logic;   	
 INT_USERCLK1_OUT    	: out std_logic;   	
 INT_USERCLK2_OUT    	: out std_logic;   	
 INT_OOBCLK_OUT      	: out std_logic;   	
 INT_MMCM_LOCK_OUT   	: out std_logic;   	
 INT_QPLLLOCK_OUT	: out std_logic_vector(1 downto 0);	
 INT_QPLLOUTCLK_OUT	: out std_logic_vector(1 downto 0);	
 INT_QPLLOUTREFCLK_OUT	: out std_logic_vector(1 downto 0);	
 INT_RXOUTCLK_OUT 	: out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	      
 INT_PCLK_SEL_SLAVE	: in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);	
     -------------Channel DRP---------------------------------
  ext_ch_gt_drpclk      : out std_logic;
  ext_ch_gt_drpaddr     : in std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*9)-1 downto 0);
  ext_ch_gt_drpen       : in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
  ext_ch_gt_drpdi       : in std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*16)-1 downto 0);
  ext_ch_gt_drpwe       : in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);

  ext_ch_gt_drpdo      : out std_logic_vector((LINK_CAP_MAX_LINK_WIDTH*16)-1 downto 0);
  ext_ch_gt_drprdy     : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);

      ---------------------------------------------------------
      -- 2. Transaction (TRN) Interface
      ---------------------------------------------------------
      -- Rx
      rx_np_ok                                 : in  std_logic;
      rx_np_req                                : in  std_logic;

      ---------------------------------------------
      -- AXI TX - RW Interface
      -----------
      s_axis_rw_tdata                          : in  std_logic_vector(C_DATA_WIDTH-1 downto 0); -- RW data from user
      s_axis_rw_tvalid                         : in  std_logic;                                 -- RW data is valid
      s_axis_rw_tready                         : out std_logic;                                 -- RW ready for data
      s_axis_rw_tstrb                          : in  std_logic_vector(STRB_WIDTH-1 downto 0);   -- RW strobe byte enables
      s_axis_rw_tlast                          : in  std_logic;                                 -- RW data is last
      s_axis_rw_tuser                          : in  std_logic_vector(3 downto 0);              -- RW user signals

      -- AXI TX - RR Interface
      -------------
      s_axis_rr_tdata                          : in  std_logic_vector(C_DATA_WIDTH-1 downto 0); -- RR data from user
      s_axis_rr_tvalid                         : in  std_logic;                                 -- RR data is valid
      s_axis_rr_tready                         : out std_logic;                                 -- RR ready for data
      s_axis_rr_tstrb                          : in  std_logic_vector(STRB_WIDTH-1 downto 0);   -- RR strobe byte enables
      s_axis_rr_tlast                          : in  std_logic;                                 -- RR data is last
      s_axis_rr_tuser                          : in  std_logic_vector(3 downto 0);              -- RR user signals

      -- AXI TX - CC Interface
      -------------
      s_axis_cc_tdata                          : in  std_logic_vector(C_DATA_WIDTH-1 downto 0); -- CC data from user
      s_axis_cc_tvalid                         : in  std_logic;                                 -- CC data is valid
      s_axis_cc_tready                         : out std_logic;                                 -- CC ready for data
      s_axis_cc_tstrb                          : in  std_logic_vector(STRB_WIDTH-1 downto 0);   -- CC strobe byte enables
      s_axis_cc_tlast                          : in  std_logic;                                 -- CC data is last
      s_axis_cc_tuser                          : in  std_logic_vector(3 downto 0);              -- CC user signals

      -- AXI RX - CW Interface
      -------------
      m_axis_cw_tdata                          : out std_logic_vector(C_DATA_WIDTH-1 downto 0); -- CW data to user
      m_axis_cw_tvalid                         : out std_logic;                                 -- CW data is valid
      m_axis_cw_tready                         : in  std_logic;                                 -- CW ready for data
      m_axis_cw_tstrb                          : out std_logic_vector(STRB_WIDTH-1 downto 0);   -- CW strobe byte enables
      m_axis_cw_tlast                          : out std_logic;                                 -- CW data is last
      m_axis_cw_tuser                          : out std_logic_vector(21 downto 0);             -- CW user signals
 
      -- AXI RX - CR Interface
      -------------
      m_axis_cr_tdata                          : out std_logic_vector(C_DATA_WIDTH-1 downto 0); -- CR data to user
      m_axis_cr_tvalid                         : out std_logic;                                 -- CR data is valid
      m_axis_cr_tready                         : in  std_logic;                                 -- CR ready for data
      m_axis_cr_tstrb                          : out std_logic_vector(STRB_WIDTH-1 downto 0);   -- CR strobe byte enables
      m_axis_cr_tlast                          : out std_logic;                                 -- CR data is last
      m_axis_cr_tuser                          : out std_logic_vector(21 downto 0);             -- CR user signals

      -- AXI RX - RC Interface
      -------------
      m_axis_rc_tdata                          : out std_logic_vector(C_DATA_WIDTH-1 downto 0); -- RC data to user
      m_axis_rc_tvalid                         : out std_logic;                                 -- RC data is valid
      m_axis_rc_tready                         : in  std_logic;                                 -- RC ready for data
      m_axis_rc_tstrb                          : out std_logic_vector(STRB_WIDTH-1 downto 0);   -- RC strobe byte enables
      m_axis_rc_tlast                          : out std_logic;                                 -- RC data is last
      m_axis_rc_tuser                          : out std_logic_vector(21 downto 0);             -- RC user signals

      -- AXI -Lite Interface - CFG Block
      ---------------------------
      s_axi_ctl_awaddr                         : in  std_logic_vector(31 downto 0);             -- AXI Lite Write address
      s_axi_ctl_awvalid                        : in  std_logic;                                 -- AXI Lite Write Address Valid
      s_axi_ctl_awready                        : out std_logic;                                 -- AXI Lite Write Address Core ready
      s_axi_ctl_wdata                          : in  std_logic_vector(31 downto 0);             -- AXI Lite Write Data
      s_axi_ctl_wstrb                          : in  std_logic_vector(3 downto 0);              -- AXI Lite Write Data strobe
      s_axi_ctl_wvalid                         : in  std_logic;                                 -- AXI Lite Write data Valid
      s_axi_ctl_wready                         : out std_logic;                                 -- AXI Lite Write Data Core ready
      s_axi_ctl_bresp                          : out std_logic_vector(1 downto 0);              -- AXI Lite Write Data strobe
      s_axi_ctl_bvalid                         : out std_logic;                                 -- AXI Lite Write data Valid
      s_axi_ctl_bready                         : in  std_logic;                                 -- AXI Lite Write Data Core ready

      s_axi_ctl_araddr                         : in  std_logic_vector(31 downto 0);             -- AXI Lite Read address
      s_axi_ctl_arvalid                        : in  std_logic;                                 -- AXI Lite Read Address Valid
      s_axi_ctl_arready                        : out std_logic;                                 -- AXI Lite Read Address Core ready
      s_axi_ctl_rdata                          : out std_logic_vector(31 downto 0);             -- AXI Lite Read Data
      s_axi_ctl_rresp                          : out std_logic_vector(1 downto 0);              -- AXI Lite Read Data strobe
      s_axi_ctl_rvalid                         : out std_logic;                                 -- AXI Lite Read data Valid
      s_axi_ctl_rready                         : in  std_logic;                                 -- AXI Lite Read Data Core ready

      -- AXI Lite User IPIC Signals
      -----------------------------
      Bus2IP_CS                                : out std_logic;                                 -- Chip Select
      Bus2IP_BE                                : out std_logic_vector(3 downto 0);              -- Byte Enable Vector
      Bus2IP_RNW                               : out std_logic;                                 -- Read Npt Write Qualifier
      Bus2IP_Addr                              : out std_logic_vector(31 downto 0);             -- Address Bus
      Bus2IP_Data                              : out std_logic_vector(31 downto 0);             -- Write Data Bus
      IP2Bus_RdAck                             : in  std_logic;                                 -- Read Acknowledgement
      IP2Bus_WrAck                             : in  std_logic;                                 -- Write Acknowledgement
      IP2Bus_Data                              : in  std_logic_vector(31 downto 0);             -- Read Data Bus
      IP2Bus_Error                             : in  std_logic;                                 -- Error Qualifier

      --Interrupts
      -------------------
      ctl_intr                                 : out std_logic;                                 -- user interrupt
      ctl_user_intr                            : in  std_logic_vector(C_NUM_USER_INTR-1 downto 0);-- User interrupt vector used only in axi_pcie_mm_s
  
      -- User Misc.
      -------------
      --user_turnoff_ok                          : in  std_logic;                                 -- Turnoff OK from user
      --user_tcfg_gnt                            : in  std_logic;                                 -- Send cfg OK from user
      np_cpl_pending                           : in  std_logic;
      RP_bridge_en                             : out std_logic;

      ---------------------------------------------------------
      -- 3. Configuration (CFG) Interface
      ---------------------------------------------------------

      blk_err_cor                              : in  std_logic;
      blk_err_ur                               : in  std_logic;
      blk_err_ecrc                             : in  std_logic;
      blk_err_cpl_timeout                      : in  std_logic;
      blk_err_cpl_abort                        : in  std_logic;
      blk_err_cpl_unexpect                     : in  std_logic;
      blk_err_posted                           : in  std_logic;
      blk_err_locked                           : in  std_logic;
      blk_err_tlp_cpl_header                   : in  std_logic_vector(47 downto 0);
      blk_err_cpl_rdy                          : out std_logic;
      blk_interrupt                            : in  std_logic;
      blk_interrupt_rdy                        : out std_logic;
      blk_interrupt_assert                     : in  std_logic;
      blk_interrupt_di                         : in  std_logic_vector(7 downto 0);
      cfg_interrupt_do                         : out std_logic_vector(7 downto 0);
      blk_interrupt_mmenable                   : out std_logic_vector(2 downto 0);
      blk_interrupt_msienable                  : out std_logic;
      blk_interrupt_msixenable                 : out std_logic;
      blk_interrupt_msixfm                     : out std_logic;
      blk_trn_pending                          : in  std_logic;
      cfg_pm_send_pme_to                       : in  std_logic;
      blk_status                               : out std_logic_vector(15 downto 0);
      blk_command                              : out std_logic_vector(15 downto 0);
      blk_dstatus                              : out std_logic_vector(15 downto 0);
      blk_dcommand                             : out std_logic_vector(15 downto 0);
      blk_lstatus                              : out std_logic_vector(15 downto 0);
      blk_lcommand                             : out std_logic_vector(15 downto 0);
      blk_dcommand2                            : out std_logic_vector(15 downto 0);
      blk_pcie_link_state                      : out std_logic_vector(2 downto 0);
      blk_dsn                                  : in  std_logic_vector(63 downto 0);
      blk_pmcsr_pme_en                         : out std_logic;
      blk_pmcsr_pme_status                     : out std_logic;
      blk_pmcsr_powerstate                     : out std_logic_vector(1 downto 0);

      cfg_msg_received                         : out std_logic;
      blk_msg_data                             : out std_logic_vector(15 downto 0);
      blk_msg_received_err_cor                 : out std_logic;
      blk_msg_received_err_non_fatal           : out std_logic;
      blk_msg_received_err_fatal               : out std_logic;
      blk_msg_received_pme_to_ack              : out std_logic;
      blk_msg_received_assert_inta             : out std_logic;
      blk_msg_received_assert_intb             : out std_logic;
      blk_msg_received_assert_intc             : out std_logic;
      blk_msg_received_assert_intd             : out std_logic;
      blk_msg_received_deassert_inta           : out std_logic;
      blk_msg_received_deassert_intb           : out std_logic;
      blk_msg_received_deassert_intc           : out std_logic;
      blk_msg_received_deassert_intd           : out std_logic;

      blk_link_up                              : out std_logic;

      blk_ds_bus_number                        : in  std_logic_vector(7 downto 0);
      blk_ds_device_number                     : in  std_logic_vector(4 downto 0);

      -- Only for End point Cores
      blk_to_turnoff                           : out  std_logic;
      blk_turnoff_ok                           : in std_logic;
      blk_pm_wake                              : in std_logic;

      blk_bus_number                           : out std_logic_vector(7 downto 0);
      blk_device_number                        : out std_logic_vector(4 downto 0);
      blk_function_number                      : out std_logic_vector(2 downto 0);

      ---------------------------------------------------------
      -- 4. Physical Layer Control and Status (PL) Interface
      ---------------------------------------------------------

      blk_pl_initial_link_width                : out std_logic_vector(2 downto 0);
      blk_pl_lane_reversal_mode                : out std_logic_vector(1 downto 0);
      blk_pl_link_gen2_capable                 : out std_logic;
      blk_pl_link_partner_gen2_supported       : out std_logic;
      blk_pl_link_upcfg_capable                : out std_logic;
      blk_pl_ltssm_state                       : out std_logic_vector(5 downto 0);
      blk_pl_sel_link_rate                     : out std_logic;
      blk_pl_sel_link_width                    : out std_logic_vector(1 downto 0);
      blk_pl_upstream_prefer_deemph            : in  std_logic;
      blk_pl_hot_rst                           : out std_logic;

      -- Flow Control
      blk_fc_cpld                              : out std_logic_vector(11 downto 0);
      blk_fc_cplh                              : out std_logic_vector(7 downto 0);
      blk_fc_npd                               : out std_logic_vector(11 downto 0);
      blk_fc_nph                               : out std_logic_vector(7 downto 0);
      blk_fc_pd                                : out std_logic_vector(11 downto 0);
      blk_fc_ph                                : out std_logic_vector(7 downto 0);
      blk_fc_sel                               : in  std_logic_vector(2 downto 0);

      -- Tx

      blk_tbuf_av                              : out std_logic_vector(5 downto 0);
      blk_tcfg_req                             : out std_logic;                                    
      blk_tcfg_gnt                             : in  std_logic;                               

      tx_err_drop                              : out std_logic;                     

      --S-6 Specific

      cfg_do                                   : out std_logic_vector(31 downto 0);
      cfg_rd_wr_done                           : out std_logic;                                
      cfg_dwaddr                               : in  std_logic_vector(9 downto 0);
      cfg_rd_en                                : in  std_logic;                          

      ---------------------------------------------------------
      -- 5. System  (SYS) Interface
      ---------------------------------------------------------

      com_sysclk                               : in  std_logic;
      com_sysrst                               : in  std_logic;
      mmcm_lock                                : out std_logic;
      com_iclk                                 : out std_logic;
      com_cclk                                 : out std_logic;
      com_corereset                            : out std_logic;

      ---------------------------------------------------------
      -- 6. Additional Signals for K7
      ---------------------------------------------------------

      clk_fab_refclk                           : in std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      clk_pclk                                 : in std_logic;
      clk_rxusrclk                             : in std_logic;
      clk_dclk                                 : in std_logic;
      clk_userclk1                             : in std_logic;
      clk_userclk2                             : in std_logic;
      clk_oobclk_in                            : in std_logic;
      clk_mmcm_lock                            : in std_logic;
      clk_txoutclk                             : out std_logic;
      clk_rxoutclk                             : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      clk_pclk_sel                             : out std_logic_vector(LINK_CAP_MAX_LINK_WIDTH-1 downto 0);
      clk_gen3                                 : out std_logic;
      PIPE_MMCM_RST_N                          : in std_logic;
      user_clk_out                             : out std_logic;
      user_reset_out                           : out std_logic;
      cfg_received_func_lvl_rst                : out std_logic;
      cfg_err_atomic_egress_blocked            : in std_logic;
      cfg_err_internal_cor                     : in std_logic;
      cfg_err_malformed                        : in std_logic;
      cfg_err_mc_blocked                       : in std_logic;
      cfg_err_poisoned                         : in std_logic;
      cfg_err_norecovery                       : in std_logic;
      cfg_err_acs                              : in std_logic;
      cfg_err_internal_uncor                   : in std_logic;
      cfg_pm_halt_aspm_l0s                     : in std_logic;
      cfg_pm_halt_aspm_l1                      : in std_logic;
      cfg_pm_force_state_en                    : in std_logic;
      cfg_pm_force_state                       : in std_logic_vector(1 downto 0);
      cfg_interrupt_stat                       : in std_logic;
      cfg_pciecap_interrupt_msgnum             : in std_logic_vector(4 downto 0);
      cfg_bridge_serr_en                       : out std_logic;
      cfg_slot_control_electromech_il_ctl_pulse: out std_logic;
      cfg_root_control_syserr_corr_err_en      : out std_logic;
      cfg_root_control_syserr_non_fatal_err_en : out std_logic;
      cfg_root_control_syserr_fatal_err_en     : out std_logic;
      cfg_root_control_pme_int_en              : out std_logic;
      cfg_aer_rooterr_corr_err_reporting_en    : out std_logic;
      cfg_aer_rooterr_non_fatal_err_reporting_en : out std_logic;
      cfg_aer_rooterr_fatal_err_reporting_en   : out std_logic;
      cfg_aer_rooterr_corr_err_received        : out std_logic;
      cfg_aer_rooterr_non_fatal_err_received   : out std_logic;
      cfg_aer_rooterr_fatal_err_received       : out std_logic;
      cfg_msg_received_pm_as_nak               : out std_logic;
      cfg_msg_received_pm_pme                  : out std_logic;
      cfg_msg_received_setslotpowerlimit       : out std_logic;
      pl_phy_lnk_up                            : out std_logic;
      pl_tx_pm_state                           : out std_logic_vector(2 downto 0);
      pl_rx_pm_state                           : out std_logic_vector(1 downto 0);
      pl_directed_change_done                  : out std_logic;
      pl_downstream_deemph_source              : in std_logic;
      cfg_err_aer_headerlog                    : in std_logic_vector(127 downto 0);
      cfg_aer_interrupt_msgnum                 : in std_logic_vector(4 downto 0);
      cfg_err_aer_headerlog_set                : out std_logic;
      cfg_aer_ecrc_check_en                    : out std_logic;
      cfg_aer_ecrc_gen_en                      : out std_logic;
      cfg_vc_tcvc_map                          : out std_logic_vector(6 downto 0);
      config_gen_req                           : out std_logic
   );
end component;

begin

   comp_enhanced_core_top_wrap : axi_pcie_v2_9_14_enhanced_core_top_wrap
      generic map (
      C_DATA_WIDTH                             => C_DATA_WIDTH,
      STRB_WIDTH                               => STRB_WIDTH,
      BAR0_U                                   => BAR0_U,
      BAR0_L                                   => BAR0_L,
      BAR1_U                                   => BAR1_U,
      BAR1_L                                   => BAR1_L,
      BAR2_U                                   => BAR2_U,
      BAR2_L                                   => BAR2_L,
      BAR3_U                                   => BAR3_U,
      BAR3_L                                   => BAR3_L,
      BAR4_U                                   => BAR4_U,
      BAR4_L                                   => BAR4_L,
      BAR5_U                                   => BAR5_U,
      BAR5_L                                   => BAR5_L,

      CARDBUS_CIS_POINTER                      => CARDBUS_CIS_POINTER,
      CLASS_CODE                               => CLASS_CODE,
      CMD_INTX_IMPLEMENTED                     => CMD_INTX_IMPLEMENTED,
      CPL_TIMEOUT_DISABLE_SUPPORTED            => CPL_TIMEOUT_DISABLE_SUPPORTED,
      CPL_TIMEOUT_RANGES_SUPPORTED             => CPL_TIMEOUT_RANGES_SUPPORTED,

      DEV_CAP_EXT_TAG_SUPPORTED                => DEV_CAP_EXT_TAG_SUPPORTED,
      DEV_CAP_MAX_PAYLOAD_SUPPORTED            => DEV_CAP_MAX_PAYLOAD_SUPPORTED,
      DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT        => DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT,
      DEVICE_ID                                => DEVICE_ID,

      DISABLE_LANE_REVERSAL                    => DISABLE_LANE_REVERSAL,
      DISABLE_SCRAMBLING                       => DISABLE_SCRAMBLING,
      DSN_BASE_PTR                             => DSN_BASE_PTR,
      DSN_CAP_NEXTPTR                          => DSN_CAP_NEXTPTR,
      DSN_CAP_ON                               => DSN_CAP_ON,

      ENABLE_MSG_ROUTE                         => ENABLE_MSG_ROUTE,
      ENABLE_RX_TD_ECRC_TRIM                   => ENABLE_RX_TD_ECRC_TRIM,
      EXPANSION_ROM_U                          => EXPANSION_ROM_U,
      EXPANSION_ROM_L                          => EXPANSION_ROM_L,
      EXT_CFG_CAP_PTR                          => EXT_CFG_CAP_PTR,
      EXT_CFG_XP_CAP_PTR                       => EXT_CFG_XP_CAP_PTR,
      HEADER_TYPE                              => HEADER_TYPE,
      INTERRUPT_PIN                            => INTERRUPT_PIN,

      LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP   => LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP,
      LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP => LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP,
      LINK_CAP_MAX_LINK_SPEED                  => LINK_CAP_MAX_LINK_SPEED,
      LINK_CAP_MAX_LINK_WIDTH                  => LINK_CAP_MAX_LINK_WIDTH,
      LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE     => LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE,

      LINK_CONTROL_RCB                         => LINK_CONTROL_RCB,
      LINK_CTRL2_DEEMPHASIS                    => LINK_CTRL2_DEEMPHASIS,
      LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE   => LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE,
      LINK_CTRL2_TARGET_LINK_SPEED             => LINK_CTRL2_TARGET_LINK_SPEED,
      LINK_STATUS_SLOT_CLOCK_CONFIG            => LINK_STATUS_SLOT_CLOCK_CONFIG,

      LL_ACK_TIMEOUT                           => LL_ACK_TIMEOUT,
      LL_ACK_TIMEOUT_EN                        => LL_ACK_TIMEOUT_EN,
      LL_ACK_TIMEOUT_FUNC                      => LL_ACK_TIMEOUT_FUNC,
      LL_REPLAY_TIMEOUT                        => LL_REPLAY_TIMEOUT,
      LL_REPLAY_TIMEOUT_EN                     => LL_REPLAY_TIMEOUT_EN,
      LL_REPLAY_TIMEOUT_FUNC                   => LL_REPLAY_TIMEOUT_FUNC,

      LTSSM_MAX_LINK_WIDTH                     => LTSSM_MAX_LINK_WIDTH,
      MSI_DECODE_ENABLE                        => MSI_DECODE_ENABLE,
      MSI_CAP_MULTIMSGCAP                      => MSI_CAP_MULTIMSGCAP,
      MSI_CAP_MULTIMSG_EXTENSION               => MSI_CAP_MULTIMSG_EXTENSION,
      MSI_CAP_ON                               => MSI_CAP_ON,
      MSI_CAP_PER_VECTOR_MASKING_CAPABLE       => MSI_CAP_PER_VECTOR_MASKING_CAPABLE,
      MSI_CAP_64_BIT_ADDR_CAPABLE              => MSI_CAP_64_BIT_ADDR_CAPABLE,

      MSIX_CAP_ON                              => MSIX_CAP_ON,
      MSIX_CAP_PBA_BIR                         => MSIX_CAP_PBA_BIR,
      MSIX_CAP_PBA_OFFSET                      => MSIX_CAP_PBA_OFFSET,
      MSIX_CAP_TABLE_BIR                       => MSIX_CAP_TABLE_BIR,
      MSIX_CAP_TABLE_OFFSET                    => MSIX_CAP_TABLE_OFFSET,
      MSIX_CAP_TABLE_SIZE                      => MSIX_CAP_TABLE_SIZE,

      PCIE_CAP_DEVICE_PORT_TYPE                => PCIE_CAP_DEVICE_PORT_TYPE,
      PCIE_CAP_INT_MSG_NUM                     => PCIE_CAP_INT_MSG_NUM,
      PCIE_CAP_NEXTPTR                         => PCIE_CAP_NEXTPTR,
      PCIE_DRP_ENABLE                          => PCIE_DRP_ENABLE,
      PIPE_PIPELINE_STAGES                     => PIPE_PIPELINE_STAGES,

      PM_CAP_DSI                               => PM_CAP_DSI,
      PM_CAP_D1SUPPORT                         => PM_CAP_D1SUPPORT,
      PM_CAP_D2SUPPORT                         => PM_CAP_D2SUPPORT,
      PM_CAP_NEXTPTR                           => PM_CAP_NEXTPTR,
      PM_CAP_PMESUPPORT                        => PM_CAP_PMESUPPORT,
      PM_CSR_NOSOFTRST                         => PM_CSR_NOSOFTRST,

      PM_DATA_SCALE0                           => PM_DATA_SCALE0,
      PM_DATA_SCALE1                           => PM_DATA_SCALE1,
      PM_DATA_SCALE2                           => PM_DATA_SCALE2,
      PM_DATA_SCALE3                           => PM_DATA_SCALE3,
      PM_DATA_SCALE4                           => PM_DATA_SCALE4,
      PM_DATA_SCALE5                           => PM_DATA_SCALE5,
      PM_DATA_SCALE6                           => PM_DATA_SCALE6,
      PM_DATA_SCALE7                           => PM_DATA_SCALE7,

      PM_DATA0                                 => PM_DATA0,
      PM_DATA1                                 => PM_DATA1,
      PM_DATA2                                 => PM_DATA2,
      PM_DATA3                                 => PM_DATA3,
      PM_DATA4                                 => PM_DATA4,
      PM_DATA5                                 => PM_DATA5,
      PM_DATA6                                 => PM_DATA6,
      PM_DATA7                                 => PM_DATA7,

      REF_CLK_FREQ                             => REF_CLK_FREQ,
      REVISION_ID                              => REVISION_ID,
      ROOT_CAP_CRS_SW_VISIBILITY               => ROOT_CAP_CRS_SW_VISIBILITY,
      SPARE_BIT0                               => SPARE_BIT0,
      SUBSYSTEM_ID                             => SUBSYSTEM_ID,
      SUBSYSTEM_VENDOR_ID                      => SUBSYSTEM_VENDOR_ID,

      SLOT_CAP_ATT_BUTTON_PRESENT              => SLOT_CAP_ATT_BUTTON_PRESENT,
      SLOT_CAP_ATT_INDICATOR_PRESENT           => SLOT_CAP_ATT_INDICATOR_PRESENT,
      SLOT_CAP_ELEC_INTERLOCK_PRESENT          => SLOT_CAP_ELEC_INTERLOCK_PRESENT,
      SLOT_CAP_HOTPLUG_CAPABLE                 => SLOT_CAP_HOTPLUG_CAPABLE,
      SLOT_CAP_HOTPLUG_SURPRISE                => SLOT_CAP_HOTPLUG_SURPRISE,
      SLOT_CAP_MRL_SENSOR_PRESENT              => SLOT_CAP_MRL_SENSOR_PRESENT,
      SLOT_CAP_NO_CMD_COMPLETED_SUPPORT        => SLOT_CAP_NO_CMD_COMPLETED_SUPPORT,
      SLOT_CAP_PHYSICAL_SLOT_NUM               => SLOT_CAP_PHYSICAL_SLOT_NUM,
      SLOT_CAP_POWER_CONTROLLER_PRESENT        => SLOT_CAP_POWER_CONTROLLER_PRESENT,
      SLOT_CAP_POWER_INDICATOR_PRESENT         => SLOT_CAP_POWER_INDICATOR_PRESENT,
      SLOT_CAP_SLOT_POWER_LIMIT_SCALE          => SLOT_CAP_SLOT_POWER_LIMIT_SCALE,
      SLOT_CAP_SLOT_POWER_LIMIT_VALUE          => SLOT_CAP_SLOT_POWER_LIMIT_VALUE,

      TL_RX_RAM_RADDR_LATENCY                  => TL_RX_RAM_RADDR_LATENCY,
      TL_RX_RAM_RDATA_LATENCY                  => TL_RX_RAM_RDATA_LATENCY,
      TL_RX_RAM_WRITE_LATENCY                  => TL_RX_RAM_WRITE_LATENCY,
      TL_TX_RAM_RADDR_LATENCY                  => TL_TX_RAM_RADDR_LATENCY,
      TL_TX_RAM_RDATA_LATENCY                  => TL_TX_RAM_RDATA_LATENCY,
      TL_TX_RAM_WRITE_LATENCY                  => TL_TX_RAM_WRITE_LATENCY,

      UPCONFIG_CAPABLE                         => UPCONFIG_CAPABLE,
      UPSTREAM_FACING                          => UPSTREAM_FACING,
      USER_CLK_FREQ                            => USER_CLK_FREQ,
      VC_BASE_PTR                              => VC_BASE_PTR,
      VC_CAP_NEXTPTR                           => VC_CAP_NEXTPTR,
      VC_CAP_ON                                => VC_CAP_ON,
      VC_CAP_REJECT_SNOOP_TRANSACTIONS         => VC_CAP_REJECT_SNOOP_TRANSACTIONS,

      VC0_CPL_INFINITE                         => VC0_CPL_INFINITE,
      VC0_RX_RAM_LIMIT                         => VC0_RX_RAM_LIMIT,
      VC0_TOTAL_CREDITS_CD                     => VC0_TOTAL_CREDITS_CD,
      VC0_TOTAL_CREDITS_CH                     => VC0_TOTAL_CREDITS_CH,
      VC0_TOTAL_CREDITS_NPH                    => VC0_TOTAL_CREDITS_NPH,
      VC0_TOTAL_CREDITS_PD                     => VC0_TOTAL_CREDITS_PD,
      VC0_TOTAL_CREDITS_PH                     => VC0_TOTAL_CREDITS_PH,
      VC0_TX_LASTPACKET                        => VC0_TX_LASTPACKET,

      VENDOR_ID                                => VENDOR_ID,
      VSEC_BASE_PTR                            => VSEC_BASE_PTR,
      VSEC_CAP_NEXTPTR                         => VSEC_CAP_NEXTPTR,
      VSEC_CAP_ON                              => VSEC_CAP_ON,

      ALLOW_X8_GEN2                            => ALLOW_X8_GEN2,
      AER_BASE_PTR                             => AER_BASE_PTR,
      AER_CAP_ECRC_CHECK_CAPABLE               => AER_CAP_ECRC_CHECK_CAPABLE,
      AER_CAP_ECRC_GEN_CAPABLE                 => AER_CAP_ECRC_GEN_CAPABLE,
      AER_CAP_ID                               => AER_CAP_ID,
      AER_CAP_INT_MSG_NUM_MSI                  => AER_CAP_INT_MSG_NUM_MSI,
      AER_CAP_INT_MSG_NUM_MSIX                 => AER_CAP_INT_MSG_NUM_MSIX,
      AER_CAP_NEXTPTR                          => AER_CAP_NEXTPTR,
      AER_CAP_ON                               => AER_CAP_ON,
      AER_CAP_PERMIT_ROOTERR_UPDATE            => AER_CAP_PERMIT_ROOTERR_UPDATE,
      AER_CAP_VERSION                          => AER_CAP_VERSION,

      CAPABILITIES_PTR                         => CAPABILITIES_PTR,
      CRM_MODULE_RSTS                          => CRM_MODULE_RSTS,
      DEV_CAP_ENDPOINT_L0S_LATENCY             => DEV_CAP_ENDPOINT_L0S_LATENCY,
      DEV_CAP_ENDPOINT_L1_LATENCY              => DEV_CAP_ENDPOINT_L1_LATENCY,
      DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE     => DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE,
      DEV_CAP_ROLE_BASED_ERROR                 => DEV_CAP_ROLE_BASED_ERROR,
      DEV_CAP_RSVD_14_12                       => DEV_CAP_RSVD_14_12,
      DEV_CAP_RSVD_17_16                       => DEV_CAP_RSVD_17_16,
      DEV_CAP_RSVD_31_29                       => DEV_CAP_RSVD_31_29,
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE      => DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE,
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE      => DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE,
      DEV_CONTROL_AUX_POWER_SUPPORTED          => DEV_CONTROL_AUX_POWER_SUPPORTED,

      DISABLE_ASPM_L1_TIMER                    => DISABLE_ASPM_L1_TIMER,
      DISABLE_BAR_FILTERING                    => DISABLE_BAR_FILTERING,
      DISABLE_ID_CHECK                         => DISABLE_ID_CHECK,
      DISABLE_RX_TC_FILTER                     => DISABLE_RX_TC_FILTER,
      DNSTREAM_LINK_NUM                        => DNSTREAM_LINK_NUM,

      DS_PORT_HOT_RST                          => DS_PORT_HOT_RST,
      DSN_CAP_ID                               => DSN_CAP_ID,
      DSN_CAP_VERSION                          => DSN_CAP_VERSION,
      ENTER_RVRY_EI_L0                         => ENTER_RVRY_EI_L0,
      INFER_EI                                 => INFER_EI,
      IS_SWITCH                                => IS_SWITCH,

      LAST_CONFIG_DWORD                        => LAST_CONFIG_DWORD,
      LINK_CAP_ASPM_SUPPORT                    => LINK_CAP_ASPM_SUPPORT,
      LINK_CAP_CLOCK_POWER_MANAGEMENT          => LINK_CAP_CLOCK_POWER_MANAGEMENT,
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    => LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1,
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    => LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2,
      LINK_CAP_L0S_EXIT_LATENCY_GEN1           => LINK_CAP_L0S_EXIT_LATENCY_GEN1,
      LINK_CAP_L0S_EXIT_LATENCY_GEN2           => LINK_CAP_L0S_EXIT_LATENCY_GEN2,
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1     => LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1,
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2     => LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2,
      LINK_CAP_L1_EXIT_LATENCY_GEN1            => LINK_CAP_L1_EXIT_LATENCY_GEN1,
      LINK_CAP_L1_EXIT_LATENCY_GEN2            => LINK_CAP_L1_EXIT_LATENCY_GEN2,
      LINK_CAP_RSVD_23_22                      => LINK_CAP_RSVD_23_22,

      MSI_BASE_PTR                             => MSI_BASE_PTR,
      MSI_CAP_ID                               => MSI_CAP_ID,
      MSI_CAP_NEXTPTR                          => MSI_CAP_NEXTPTR,
      MSIX_BASE_PTR                            => MSIX_BASE_PTR,
      MSIX_CAP_ID                              => MSIX_CAP_ID,
      MSIX_CAP_NEXTPTR                         => MSIX_CAP_NEXTPTR,
      N_FTS_COMCLK_GEN1                        => N_FTS_COMCLK_GEN1,
      N_FTS_COMCLK_GEN2                        => N_FTS_COMCLK_GEN2,
      N_FTS_GEN1                               => N_FTS_GEN1,
      N_FTS_GEN2                               => N_FTS_GEN2,

      PCIE_BASE_PTR                            => PCIE_BASE_PTR,
      PCIE_CAP_CAPABILITY_ID                   => PCIE_CAP_CAPABILITY_ID,
      PCIE_CAP_CAPABILITY_VERSION              => PCIE_CAP_CAPABILITY_VERSION,
      PCIE_CAP_ON                              => PCIE_CAP_ON,
      PCIE_CAP_RSVD_15_14                      => PCIE_CAP_RSVD_15_14,
      PCIE_CAP_SLOT_IMPLEMENTED                => PCIE_CAP_SLOT_IMPLEMENTED,
      PCIE_REVISION                            => PCIE_REVISION,
      PGL0_LANE                                => PGL0_LANE,
      PGL1_LANE                                => PGL1_LANE,
      PGL2_LANE                                => PGL2_LANE,
      PGL3_LANE                                => PGL3_LANE,
      PGL4_LANE                                => PGL4_LANE,
      PGL5_LANE                                => PGL5_LANE,
      PGL6_LANE                                => PGL6_LANE,
      PGL7_LANE                                => PGL7_LANE,
      PL_AUTO_CONFIG                           => PL_AUTO_CONFIG,
      PL_FAST_TRAIN                            => PL_FAST_TRAIN,
      PCIE_EXT_CLK                             => PCIE_EXT_CLK,
       PCIE_EXT_GT_COMMON     =>PCIE_EXT_GT_COMMON ,
       EXT_CH_GT_DRP            => EXT_CH_GT_DRP,	    
      NO_SLV_ERR                               => NO_SLV_ERR,

 TX_MARGIN_FULL_0  =>TX_MARGIN_FULL_0  ,
 TX_MARGIN_FULL_1  =>TX_MARGIN_FULL_1  ,
 TX_MARGIN_FULL_2  =>TX_MARGIN_FULL_2  ,
 TX_MARGIN_FULL_3  =>TX_MARGIN_FULL_3  ,
 TX_MARGIN_FULL_4  =>TX_MARGIN_FULL_4  ,
 TX_MARGIN_LOW_0   =>TX_MARGIN_LOW_0   ,
 TX_MARGIN_LOW_1   =>TX_MARGIN_LOW_1   ,
 TX_MARGIN_LOW_2   =>TX_MARGIN_LOW_2   ,
 TX_MARGIN_LOW_3   =>TX_MARGIN_LOW_3   ,
 TX_MARGIN_LOW_4   =>TX_MARGIN_LOW_4   ,
      PM_BASE_PTR                              => PM_BASE_PTR,
      PM_CAP_AUXCURRENT                        => PM_CAP_AUXCURRENT,
      PM_CAP_ID                                => PM_CAP_ID,
      PM_CAP_ON                                => PM_CAP_ON,
      PM_CAP_PME_CLOCK                         => PM_CAP_PME_CLOCK,
      PM_CAP_RSVD_04                           => PM_CAP_RSVD_04,
      PM_CAP_VERSION                           => PM_CAP_VERSION,
      PM_CSR_BPCCEN                            => PM_CSR_BPCCEN,
      PM_CSR_B2B3                              => PM_CSR_B2B3,

      RECRC_CHK                                => RECRC_CHK,
      RECRC_CHK_TRIM                           => RECRC_CHK_TRIM,
      SELECT_DLL_IF                            => SELECT_DLL_IF,
      SPARE_BIT1                               => SPARE_BIT1,
      SPARE_BIT2                               => SPARE_BIT2,
      SPARE_BIT3                               => SPARE_BIT3,
      SPARE_BIT4                               => SPARE_BIT4,
      SPARE_BIT5                               => SPARE_BIT5,
      SPARE_BIT6                               => SPARE_BIT6,
      SPARE_BIT7                               => SPARE_BIT7,
      SPARE_BIT8                               => SPARE_BIT8,
      SPARE_BYTE0                              => SPARE_BYTE0,
      SPARE_BYTE1                              => SPARE_BYTE1,
      SPARE_BYTE2                              => SPARE_BYTE2,
      SPARE_BYTE3                              => SPARE_BYTE3,
      SPARE_WORD0                              => SPARE_WORD0,
      SPARE_WORD1                              => SPARE_WORD1,
      SPARE_WORD2                              => SPARE_WORD2,
      SPARE_WORD3                              => SPARE_WORD3,

      TL_RBYPASS                               => TL_RBYPASS,
      TL_TFC_DISABLE                           => TL_TFC_DISABLE,
      TL_TX_CHECKS_DISABLE                     => TL_TX_CHECKS_DISABLE,
      EXIT_LOOPBACK_ON_EI                      => EXIT_LOOPBACK_ON_EI,
      UR_INV_REQ                               => UR_INV_REQ,

      VC_CAP_ID                                => VC_CAP_ID,
      VC_CAP_VERSION                           => VC_CAP_VERSION,
      VSEC_CAP_HDR_ID                          => VSEC_CAP_HDR_ID,
      VSEC_CAP_HDR_LENGTH                      => VSEC_CAP_HDR_LENGTH,
      VSEC_CAP_HDR_REVISION                    => VSEC_CAP_HDR_REVISION,
      VSEC_CAP_ID                              => VSEC_CAP_ID,
      VSEC_CAP_IS_LINK_VISIBLE                 => VSEC_CAP_IS_LINK_VISIBLE,
      VSEC_CAP_VERSION                         => VSEC_CAP_VERSION,

      C_BASEADDR_U                             => C_BASEADDR_U,
      C_BASEADDR_L                             => C_BASEADDR_L,
      C_HIGHADDR_U                             => C_HIGHADDR_U,
      C_HIGHADDR_L                             => C_HIGHADDR_L,

      C_MAX_LNK_WDT                            => C_MAX_LNK_WDT,
      C_ROOT_PORT                              => C_ROOT_PORT,
      C_RP_BAR_HIDE                            => C_RP_BAR_HIDE,
      C_RX_REALIGN                             => C_RX_REALIGN,
      C_RX_PRESERVE_ORDER                      => C_RX_PRESERVE_ORDER,
      C_LAST_CORE_CAP_ADDR                     => C_LAST_CORE_CAP_ADDR,
      C_VSEC_CAP_ADDR                          => C_VSEC_CAP_ADDR,
      C_VSEC_CAP_LAST                          => C_VSEC_CAP_LAST,
      C_VSEC_ID                                => C_VSEC_ID,
      C_DEVICE_NUMBER                          => C_DEVICE_NUMBER,
      C_NUM_USER_INTR                          => C_NUM_USER_INTR,
      C_USER_PTR                               => C_USER_PTR,
      C_COMP_TIMEOUT                           => C_COMP_TIMEOUT,
      PTR_WIDTH                                => PTR_WIDTH,
      C_FAMILY                                 => C_FAMILY,

      USR_CFG                                  => USR_CFG,
      USR_EXT_CFG                              => USR_EXT_CFG,
      LINK_CAP_L0S_EXIT_LATENCY                => LINK_CAP_L0S_EXIT_LATENCY,
      LINK_CAP_L1_EXIT_LATENCY                 => LINK_CAP_L1_EXIT_LATENCY,
      PLM_AUTO_CONFIG                          => PLM_AUTO_CONFIG,
      FAST_TRAIN                               => FAST_TRAIN,
      PCIE_GENERIC                             => PCIE_GENERIC,
      GTP_SEL                                  => GTP_SEL,
      CFG_VEN_ID                               => CFG_VEN_ID,
      CFG_DEV_ID                               => CFG_DEV_ID,
      CFG_REV_ID                               => CFG_REV_ID,
      CFG_SUBSYS_VEN_ID                        => CFG_SUBSYS_VEN_ID,
      CFG_SUBSYS_ID                            => CFG_SUBSYS_ID,

      AER_CAP_MULTIHEADER                      => AER_CAP_MULTIHEADER,
      AER_CAP_OPTIONAL_ERR_SUPPORT             => AER_CAP_OPTIONAL_ERR_SUPPORT,
      DEV_CAP2_ARI_FORWARDING_SUPPORTED        => DEV_CAP2_ARI_FORWARDING_SUPPORTED,
      DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED  => DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED,
      DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED  => DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED,
      DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED      => DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED,
      DEV_CAP2_CAS128_COMPLETER_SUPPORTED      => DEV_CAP2_CAS128_COMPLETER_SUPPORTED,
      DEV_CAP2_TPH_COMPLETER_SUPPORTED         => DEV_CAP2_TPH_COMPLETER_SUPPORTED,
      DEV_CONTROL_EXT_TAG_DEFAULT              => DEV_CONTROL_EXT_TAG_DEFAULT,
      DISABLE_RX_POISONED_RESP                 => DISABLE_RX_POISONED_RESP,
      LINK_CAP_ASPM_OPTIONALITY                => LINK_CAP_ASPM_OPTIONALITY,
      RBAR_BASE_PTR                            => RBAR_BASE_PTR,
      RBAR_CAP_CONTROL_ENCODEDBAR0             => RBAR_CAP_CONTROL_ENCODEDBAR0,
      RBAR_CAP_CONTROL_ENCODEDBAR1             => RBAR_CAP_CONTROL_ENCODEDBAR1,
      RBAR_CAP_CONTROL_ENCODEDBAR2             => RBAR_CAP_CONTROL_ENCODEDBAR2,
      RBAR_CAP_CONTROL_ENCODEDBAR3             => RBAR_CAP_CONTROL_ENCODEDBAR3,
      RBAR_CAP_CONTROL_ENCODEDBAR4             => RBAR_CAP_CONTROL_ENCODEDBAR4,
      RBAR_CAP_CONTROL_ENCODEDBAR5             => RBAR_CAP_CONTROL_ENCODEDBAR5,
      RBAR_CAP_INDEX0                          => RBAR_CAP_INDEX0,
      RBAR_CAP_INDEX1                          => RBAR_CAP_INDEX1,
      RBAR_CAP_INDEX2                          => RBAR_CAP_INDEX2,
      RBAR_CAP_INDEX3                          => RBAR_CAP_INDEX3,
      RBAR_CAP_INDEX4                          => RBAR_CAP_INDEX4,
      RBAR_CAP_INDEX5                          => RBAR_CAP_INDEX5,
      RBAR_CAP_ON                              => RBAR_CAP_ON,
      RBAR_CAP_SUP0                            => RBAR_CAP_SUP0,
      RBAR_CAP_SUP1                            => RBAR_CAP_SUP1,
      RBAR_CAP_SUP2                            => RBAR_CAP_SUP2,
      RBAR_CAP_SUP3                            => RBAR_CAP_SUP3,
      RBAR_CAP_SUP4                            => RBAR_CAP_SUP4,
      RBAR_CAP_SUP5                            => RBAR_CAP_SUP5,
      RBAR_NUM                                 => RBAR_NUM,
      TRN_NP_FC                                => TRN_NP_FC,
      TRN_DW                                   => TRN_DW,
      UR_ATOMIC                                => UR_ATOMIC,
      UR_PRS_RESPONSE                          => UR_PRS_RESPONSE,
      USER_CLK2_DIV2                           => USER_CLK2_DIV2,
      VC0_TOTAL_CREDITS_NPD                    => VC0_TOTAL_CREDITS_NPD,
      LINK_CAP_RSVD_23                         => LINK_CAP_RSVD_23,
      CFG_ECRC_ERR_CPLSTAT                     => CFG_ECRC_ERR_CPLSTAT,
      DISABLE_ERR_MSG                          => DISABLE_ERR_MSG,
      DISABLE_LOCKED_FILTER                    => DISABLE_LOCKED_FILTER,
      DISABLE_PPM_FILTER                       => DISABLE_PPM_FILTER,
      ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED   => ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED,
      INTERRUPT_STAT_AUTO                      => INTERRUPT_STAT_AUTO,
      MPS_FORCE                                => MPS_FORCE,
      PM_ASPML0S_TIMEOUT                       => PM_ASPML0S_TIMEOUT,
      PM_ASPML0S_TIMEOUT_EN                    => PM_ASPML0S_TIMEOUT_EN,
      PM_ASPML0S_TIMEOUT_FUNC                  => PM_ASPML0S_TIMEOUT_FUNC,
      PM_ASPM_FASTEXIT                         => PM_ASPM_FASTEXIT,
      PM_MF                                    => PM_MF,
      RP_AUTO_SPD                              => RP_AUTO_SPD,
      RP_AUTO_SPD_LOOPCNT                      => RP_AUTO_SPD_LOOPCNT,
      SIM_VERSION                              => SIM_VERSION,
      SSL_MESSAGE_AUTO                         => SSL_MESSAGE_AUTO,
      TECRC_EP_INV                             => TECRC_EP_INV,
      UR_CFG1                                  => UR_CFG1,
      USE_RID_PINS                             => USE_RID_PINS,
      DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED     => DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED,
      DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED    => DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED,
      DEV_CAP2_LTR_MECHANISM_SUPPORTED         => DEV_CAP2_LTR_MECHANISM_SUPPORTED,
      DEV_CAP2_MAX_ENDEND_TLP_PREFIXES         => DEV_CAP2_MAX_ENDEND_TLP_PREFIXES,
      DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING      => DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING,
      RBAR_CAP_ID                              => RBAR_CAP_ID,
      RBAR_CAP_NEXTPTR                         => RBAR_CAP_NEXTPTR,
      RBAR_CAP_VERSION                         => RBAR_CAP_VERSION,
      PCIE_USE_MODE                            => PCIE_USE_MODE,
      PCIE_GT_DEVICE                           => PCIE_GT_DEVICE,
      PCIE_CHAN_BOND                           => PCIE_CHAN_BOND,
      PCIE_PLL_SEL                             => PCIE_PLL_SEL,
      PCIE_ASYNC_EN                            => PCIE_ASYNC_EN,
      PCIE_TXBUF_EN                            => PCIE_TXBUF_EN,
      EXT_PIPE_INTERFACE                       => EXT_PIPE_INTERFACE 
      )
      port map ( 
      -- 1. PCI Express (pci_exp) Interface
      ---------------------------------------------------------
      -- Tx
      pci_exp_txp                              => pci_exp_txp,
      pci_exp_txn                              => pci_exp_txn,
      -- Rx
      pci_exp_rxp                              => pci_exp_rxp,
      pci_exp_rxn                              => pci_exp_rxn,
 qpll_drp_crscode      => qpll_drp_crscode    ,
 qpll_drp_fsm          => qpll_drp_fsm        ,
 qpll_drp_done         => qpll_drp_done       ,
 qpll_drp_reset        => qpll_drp_reset      ,
 qpll_qplllock         => qpll_qplllock       ,
 qpll_qplloutclk       => qpll_qplloutclk     ,
 qpll_qplloutrefclk    => qpll_qplloutrefclk  ,
  qpll_qplld    => qpll_qplld    ,
  qpll_qpllreset=> qpll_qpllreset,
  qpll_drp_clk  => qpll_drp_clk  ,
  qpll_drp_rst_n=> qpll_drp_rst_n,
  qpll_drp_ovrd => qpll_drp_ovrd ,
  qpll_drp_gen3 => qpll_drp_gen3 ,
  qpll_drp_start=> qpll_drp_start,

  pipe_txprbssel      => pipe_txprbssel     , 
  pipe_rxprbssel      => pipe_rxprbssel     , 
  pipe_txprbsforceerr => pipe_txprbsforceerr, 
  pipe_rxprbscntreset => pipe_rxprbscntreset, 
  pipe_loopback       => pipe_loopback      , 
  pipe_txinhibit        => pipe_txinhibit       ,

  pipe_rxprbserr        => pipe_rxprbserr       ,
  pipe_rst_fsm          => pipe_rst_fsm         ,
  pipe_qrst_fsm         => pipe_qrst_fsm        ,
  pipe_rate_fsm         => pipe_rate_fsm        ,
  pipe_sync_fsm_tx      => pipe_sync_fsm_tx     ,
  pipe_sync_fsm_rx      => pipe_sync_fsm_rx     ,
  pipe_drp_fsm          => pipe_drp_fsm         ,

  pipe_rst_idle => pipe_rst_idle ,
  pipe_qrst_idle=> pipe_qrst_idle,
  pipe_rate_idle=> pipe_rate_idle,
  pipe_eyescandataerror	=> pipe_eyescandataerror,
  pipe_rxstatus    => pipe_rxstatus,
  pipe_dmonitorout => pipe_dmonitorout,
  
  pipe_cpll_lock         =>  pipe_cpll_lock 	,
  pipe_qpll_lock         =>  pipe_qpll_lock 	,
  pipe_rxpmaresetdone    =>  pipe_rxpmaresetdone	,       
  pipe_rxbufstatus 	 =>  pipe_rxbufstatus 	,         
  pipe_txphaligndone     =>  pipe_txphaligndone 	,       
  pipe_txphinitdone 	 =>  pipe_txphinitdone 	,        
  pipe_txdlysresetdone   =>  pipe_txdlysresetdone,    
  pipe_rxphaligndone     =>  pipe_rxphaligndone 	,      
  pipe_rxdlysresetdone   =>  pipe_rxdlysresetdone,     
  pipe_rxsyncdone 	 =>  pipe_rxsyncdone 	,       
  pipe_rxdisperr 	 =>  pipe_rxdisperr 	,       
  pipe_rxnotintable 	 =>  pipe_rxnotintable 	,      
  pipe_rxcommadet 	 =>  pipe_rxcommadet 	,        

  gt_ch_drp_rdy => gt_ch_drp_rdy ,
  pipe_debug_0 	=> pipe_debug_0 	,
  pipe_debug_1 	=> pipe_debug_1 	,
  pipe_debug_2 	=> pipe_debug_2 	,
  pipe_debug_3 	=> pipe_debug_3 	,
  pipe_debug_4 	=> pipe_debug_4 	,
  pipe_debug_5 	=> pipe_debug_5 	,
  pipe_debug_6 	=> pipe_debug_6 	,
  pipe_debug_7 	=> pipe_debug_7 	,
  pipe_debug_8 	=> pipe_debug_8 	,
  pipe_debug_9 	=> pipe_debug_9 	,
  pipe_debug   	=> pipe_debug   	,

  common_commands_in		=>common_commands_in	,
  pipe_rx_0_sigs		=>pipe_rx_0_sigs	,
  pipe_rx_1_sigs		=>pipe_rx_1_sigs	,
  pipe_rx_2_sigs		=>pipe_rx_2_sigs	,
  pipe_rx_3_sigs		=>pipe_rx_3_sigs	,
  pipe_rx_4_sigs		=>pipe_rx_4_sigs	,
  pipe_rx_5_sigs		=>pipe_rx_5_sigs	,
  pipe_rx_6_sigs		=>pipe_rx_6_sigs	,
  pipe_rx_7_sigs		=>pipe_rx_7_sigs	,
                                                 
  common_commands_out		=>common_commands_out	,
  pipe_tx_0_sigs		=>pipe_tx_0_sigs	,
  pipe_tx_1_sigs		=>pipe_tx_1_sigs	,
  pipe_tx_2_sigs		=>pipe_tx_2_sigs	,
  pipe_tx_3_sigs		=>pipe_tx_3_sigs	,
  pipe_tx_4_sigs		=>pipe_tx_4_sigs	,
  pipe_tx_5_sigs		=>pipe_tx_5_sigs	,
  pipe_tx_6_sigs		=>pipe_tx_6_sigs	,
  pipe_tx_7_sigs		=>pipe_tx_7_sigs	,

INT_PCLK_OUT_SLAVE	=>		INT_PCLK_OUT_SLAVE,	
INT_RXUSRCLK_OUT  	=>      	INT_RXUSRCLK_OUT  ,      
INT_RXOUTCLK_OUT  	=>      	INT_RXOUTCLK_OUT  ,      
INT_DCLK_OUT	  	=>      	INT_DCLK_OUT	  ,      
INT_USERCLK1_OUT  	=>      	INT_USERCLK1_OUT  ,      
INT_USERCLK2_OUT  	=>      	INT_USERCLK2_OUT  ,      
INT_OOBCLK_OUT	  	=>      	INT_OOBCLK_OUT	  ,      
INT_MMCM_LOCK_OUT 	=>      	INT_MMCM_LOCK_OUT ,      
INT_QPLLLOCK_OUT  	=>      	INT_QPLLLOCK_OUT  ,      
INT_QPLLOUTCLK_OUT	=>		INT_QPLLOUTCLK_OUT,	
INT_QPLLOUTREFCLK_OUT		=>	INT_QPLLOUTREFCLK_OUT,	
INT_PCLK_SEL_SLAVE		=>	INT_PCLK_SEL_SLAVE   ,   

     -------------Channel DRP---------------------------------
  ext_ch_gt_drpclk    => ext_ch_gt_drpclk ,
  ext_ch_gt_drpaddr   => ext_ch_gt_drpaddr,
  ext_ch_gt_drpen     => ext_ch_gt_drpen  ,
  ext_ch_gt_drpdi     => ext_ch_gt_drpdi  ,
  ext_ch_gt_drpwe     => ext_ch_gt_drpwe  ,
                                          
  ext_ch_gt_drpdo     => ext_ch_gt_drpdo  ,
  ext_ch_gt_drprdy    => ext_ch_gt_drprdy ,

      ---------------------------------------------------------
      -- 2. Transaction (TRN) Interface
      ---------------------------------------------------------
      -- Rx
      rx_np_ok                                 => rx_np_ok,
      rx_np_req                                => rx_np_req,

      ---------------------------------------------
      -- AXI TX - RW Interface
      -----------
      s_axis_rw_tdata                          => s_axis_rw_tdata,
      s_axis_rw_tvalid                         => s_axis_rw_tvalid,
      s_axis_rw_tready                         => s_axis_rw_tready,
      s_axis_rw_tstrb                          => s_axis_rw_tstrb,
      s_axis_rw_tlast                          => s_axis_rw_tlast,
      s_axis_rw_tuser                          => s_axis_rw_tuser,

      -- AXI TX - RR Interface
      -------------
      s_axis_rr_tdata                          => s_axis_rr_tdata,
      s_axis_rr_tvalid                         => s_axis_rr_tvalid,
      s_axis_rr_tready                         => s_axis_rr_tready,
      s_axis_rr_tstrb                          => s_axis_rr_tstrb,
      s_axis_rr_tlast                          => s_axis_rr_tlast,
      s_axis_rr_tuser                          => s_axis_rr_tuser,

      -- AXI TX - CC Interface
      -------------
      s_axis_cc_tdata                          => s_axis_cc_tdata,
      s_axis_cc_tvalid                         => s_axis_cc_tvalid,
      s_axis_cc_tready                         => s_axis_cc_tready,
      s_axis_cc_tstrb                          => s_axis_cc_tstrb,
      s_axis_cc_tlast                          => s_axis_cc_tlast,
      s_axis_cc_tuser                          => s_axis_cc_tuser,

      -- AXI RX - CW Interface
      -------------
      m_axis_cw_tdata                          => m_axis_cw_tdata,
      m_axis_cw_tvalid                         => m_axis_cw_tvalid,
      m_axis_cw_tready                         => m_axis_cw_tready,
      m_axis_cw_tstrb                          => m_axis_cw_tstrb,
      m_axis_cw_tlast                          => m_axis_cw_tlast,
      m_axis_cw_tuser                          => m_axis_cw_tuser,
 
      -- AXI RX - CR Interface
      -------------
      m_axis_cr_tdata                          => m_axis_cr_tdata,
      m_axis_cr_tvalid                         => m_axis_cr_tvalid,
      m_axis_cr_tready                         => m_axis_cr_tready,
      m_axis_cr_tstrb                          => m_axis_cr_tstrb,
      m_axis_cr_tlast                          => m_axis_cr_tlast,
      m_axis_cr_tuser                          => m_axis_cr_tuser,

      -- AXI RX - RC Interface
      -------------
      m_axis_rc_tdata                          => m_axis_rc_tdata,
      m_axis_rc_tvalid                         => m_axis_rc_tvalid,
      m_axis_rc_tready                         => m_axis_rc_tready,
      m_axis_rc_tstrb                          => m_axis_rc_tstrb,
      m_axis_rc_tlast                          => m_axis_rc_tlast,
      m_axis_rc_tuser                          => m_axis_rc_tuser,

      -- AXI -Lite Interface - CFG Block
      ---------------------------
      s_axi_ctl_awaddr                         => s_axi_ctl_awaddr,
      s_axi_ctl_awvalid                        => s_axi_ctl_awvalid,
      s_axi_ctl_awready                        => s_axi_ctl_awready,
      s_axi_ctl_wdata                          => s_axi_ctl_wdata,
      s_axi_ctl_wstrb                          => s_axi_ctl_wstrb,
      s_axi_ctl_wvalid                         => s_axi_ctl_wvalid,
      s_axi_ctl_wready                         => s_axi_ctl_wready,
      s_axi_ctl_bresp                          => s_axi_ctl_bresp,
      s_axi_ctl_bvalid                         => s_axi_ctl_bvalid,
      s_axi_ctl_bready                         => s_axi_ctl_bready,

      s_axi_ctl_araddr                         => s_axi_ctl_araddr,
      s_axi_ctl_arvalid                        => s_axi_ctl_arvalid,
      s_axi_ctl_arready                        => s_axi_ctl_arready,
      s_axi_ctl_rdata                          => s_axi_ctl_rdata,
      s_axi_ctl_rresp                          => s_axi_ctl_rresp,
      s_axi_ctl_rvalid                         => s_axi_ctl_rvalid,
      s_axi_ctl_rready                         => s_axi_ctl_rready,

      -- AXI Lite User IPIC Signals
      -----------------------------
      Bus2IP_CS                                => Bus2IP_CS,
      Bus2IP_BE                                => Bus2IP_BE,
      Bus2IP_RNW                               => Bus2IP_RNW,
      Bus2IP_Addr                              => Bus2IP_Addr,
      Bus2IP_Data                              => Bus2IP_Data,
      IP2Bus_RdAck                             => IP2Bus_RdAck,
      IP2Bus_WrAck                             => IP2Bus_WrAck,
      IP2Bus_Data                              => IP2Bus_Data,
      IP2Bus_Error                             => IP2Bus_Error,

      --Interrupts
      -------------------
      ctl_intr                                 => ctl_intr,
      ctl_user_intr                            => ctl_user_intr,
  
      -- User Misc.
      -------------
      --user_turnoff_ok                          => user_turnoff_ok,
      --user_tcfg_gnt                            => user_tcfg_gnt,

      np_cpl_pending                           => np_cpl_pending,
      RP_bridge_en                             => RP_bridge_en,

      ---------------------------------------------------------
      -- 3. Configuration (CFG) Interface
      ---------------------------------------------------------

      blk_err_cor                              => blk_err_cor,
      blk_err_ur                               => blk_err_ur,
      blk_err_ecrc                             => blk_err_ecrc,
      blk_err_cpl_timeout                      => blk_err_cpl_timeout,
      blk_err_cpl_abort                        => blk_err_cpl_abort,
      blk_err_cpl_unexpect                     => blk_err_cpl_unexpect,
      blk_err_posted                           => blk_err_posted,
      blk_err_locked                           => blk_err_locked,
      blk_err_tlp_cpl_header                   => blk_err_tlp_cpl_header,
      blk_err_cpl_rdy                          => blk_err_cpl_rdy,
      blk_interrupt                            => blk_interrupt,
      blk_interrupt_rdy                        => blk_interrupt_rdy,
      blk_interrupt_assert                     => blk_interrupt_assert,
      blk_interrupt_di                         => blk_interrupt_di,
      cfg_interrupt_do                         => cfg_interrupt_do,
      blk_interrupt_mmenable                   => blk_interrupt_mmenable,
      blk_interrupt_msienable                  => blk_interrupt_msienable,
      blk_interrupt_msixenable                 => blk_interrupt_msixenable,
      blk_interrupt_msixfm                     => blk_interrupt_msixfm,
      blk_trn_pending                          => blk_trn_pending,
      cfg_pm_send_pme_to                       => cfg_pm_send_pme_to,
      blk_status                               => blk_status,
      blk_command                              => blk_command,
      blk_dstatus                              => blk_dstatus,
      blk_dcommand                             => blk_dcommand,
      blk_lstatus                              => blk_lstatus,
      blk_lcommand                             => blk_lcommand,
      blk_dcommand2                            => blk_dcommand2,
      blk_pcie_link_state                      => blk_pcie_link_state,
      blk_dsn                                  => blk_dsn,
      blk_pmcsr_pme_en                         => blk_pmcsr_pme_en,
      blk_pmcsr_pme_status                     => blk_pmcsr_pme_status,
      blk_pmcsr_powerstate                     => blk_pmcsr_powerstate,

      cfg_msg_received                         => cfg_msg_received,
      blk_msg_data                             => blk_msg_data,
      blk_msg_received_err_cor                 => blk_msg_received_err_cor,
      blk_msg_received_err_non_fatal           => blk_msg_received_err_non_fatal,
      blk_msg_received_err_fatal               => blk_msg_received_err_fatal,
      blk_msg_received_pme_to_ack              => blk_msg_received_pme_to_ack,
      blk_msg_received_assert_inta             => blk_msg_received_assert_inta,
      blk_msg_received_assert_intb             => blk_msg_received_assert_intb,
      blk_msg_received_assert_intc             => blk_msg_received_assert_intc,
      blk_msg_received_assert_intd             => blk_msg_received_assert_intd,
      blk_msg_received_deassert_inta           => blk_msg_received_deassert_inta,
      blk_msg_received_deassert_intb           => blk_msg_received_deassert_intb,
      blk_msg_received_deassert_intc           => blk_msg_received_deassert_intc,
      blk_msg_received_deassert_intd           => blk_msg_received_deassert_intd,

      blk_link_up                              => blk_link_up,

      blk_ds_bus_number                        => blk_ds_bus_number,
      blk_ds_device_number                     => blk_ds_device_number,

      -- Only for End point Cores
      blk_to_turnoff                           => blk_to_turnoff,
      blk_turnoff_ok                           => blk_turnoff_ok,
      blk_pm_wake                              => blk_pm_wake,

      blk_bus_number                           => blk_bus_number,
      blk_device_number                        => blk_device_number,
      blk_function_number                      => blk_function_number,

      ---------------------------------------------------------
      -- 4. Physical Layer Control and Status (PL) Interface
      ---------------------------------------------------------

      blk_pl_initial_link_width                => blk_pl_initial_link_width,
      blk_pl_lane_reversal_mode                => blk_pl_lane_reversal_mode,
      blk_pl_link_gen2_capable                 => blk_pl_link_gen2_capable,
      blk_pl_link_partner_gen2_supported       => blk_pl_link_partner_gen2_supported,
      blk_pl_link_upcfg_capable                => blk_pl_link_upcfg_capable,
      blk_pl_ltssm_state                       => blk_pl_ltssm_state,
      blk_pl_sel_link_rate                     => blk_pl_sel_link_rate,
      blk_pl_sel_link_width                    => blk_pl_sel_link_width,
      blk_pl_upstream_prefer_deemph            => blk_pl_upstream_prefer_deemph,
      blk_pl_hot_rst                           => blk_pl_hot_rst,

      -- Flow Control
      blk_fc_cpld                              => blk_fc_cpld,
      blk_fc_cplh                              => blk_fc_cplh,
      blk_fc_npd                               => blk_fc_npd,
      blk_fc_nph                               => blk_fc_nph,
      blk_fc_pd                                => blk_fc_pd,
      blk_fc_ph                                => blk_fc_ph,
      blk_fc_sel                               => blk_fc_sel,

      -- Tx

      blk_tbuf_av                              => blk_tbuf_av,
      blk_tcfg_req                             => blk_tcfg_req,                 
      blk_tcfg_gnt                             => blk_tcfg_gnt,            

      tx_err_drop                              => tx_err_drop,  

      --S-6 Specific

      cfg_do                                   => cfg_do,
      cfg_rd_wr_done                           => cfg_rd_wr_done,            
      cfg_dwaddr                               => cfg_dwaddr,
      cfg_rd_en                                => cfg_rd_en,      

      ---------------------------------------------------------
      -- 5. System  (SYS) Interface
      ---------------------------------------------------------

      com_sysclk                               => com_sysclk,
      com_sysrst                               => com_sysrst,
      mmcm_lock                                => mmcm_lock,
      com_iclk                                 => com_iclk,
      com_cclk                                 => com_cclk,
      com_corereset                            => com_corereset,
      
      ---------------------------------------------------------
      -- 6. Additional Signals for K7
      ---------------------------------------------------------
      
      clk_fab_refclk                           => clk_fab_refclk,
      clk_pclk                                 => clk_pclk,
      clk_rxusrclk                             => clk_rxusrclk,
      clk_dclk                                 => clk_dclk,
      clk_userclk1                             => clk_userclk1,
      clk_userclk2                             => clk_userclk2,
      clk_oobclk_in                            => clk_oobclk_in,
      clk_mmcm_lock                            => clk_mmcm_lock,
      clk_txoutclk                             => clk_txoutclk,
      clk_rxoutclk                             => clk_rxoutclk,
      clk_pclk_sel                             => clk_pclk_sel,
      clk_gen3                                 => clk_gen3,
      PIPE_MMCM_RST_N                          => PIPE_MMCM_RST_N,
      user_clk_out                             => open,
      user_reset_out                           => open,
      cfg_received_func_lvl_rst                => open,
      cfg_err_atomic_egress_blocked            => '0',
      cfg_err_internal_cor                     => '0',
      cfg_err_malformed                        => '0',
      cfg_err_mc_blocked                       => '0',
      cfg_err_poisoned                         => '0',
      cfg_err_norecovery                       => '0',
      cfg_err_acs                              => '0',
      cfg_err_internal_uncor                   => '0',
      cfg_pm_halt_aspm_l0s                     => '0',
      cfg_pm_halt_aspm_l1                      => '0',
      cfg_pm_force_state_en                    => '0',
      cfg_pm_force_state                       => (others => '0'),
      cfg_interrupt_stat                       => '0',
      cfg_pciecap_interrupt_msgnum             => (others => '0'),
      cfg_bridge_serr_en                       => open,
      cfg_slot_control_electromech_il_ctl_pulse => open,
      cfg_root_control_syserr_corr_err_en      => open,
      cfg_root_control_syserr_non_fatal_err_en => open,
      cfg_root_control_syserr_fatal_err_en     => open,
      cfg_root_control_pme_int_en              => open,
      cfg_aer_rooterr_corr_err_reporting_en    => open,
      cfg_aer_rooterr_non_fatal_err_reporting_en => open,
      cfg_aer_rooterr_fatal_err_reporting_en   => open,
      cfg_aer_rooterr_corr_err_received        => open,
      cfg_aer_rooterr_non_fatal_err_received   => open,
      cfg_aer_rooterr_fatal_err_received       => open,
      cfg_msg_received_pm_as_nak               => open,
      cfg_msg_received_pm_pme                  => open,
      cfg_msg_received_setslotpowerlimit       => open,
      pl_phy_lnk_up                            => open,
      pl_tx_pm_state                           => open,
      pl_rx_pm_state                           => open,
      pl_directed_change_done                  => open,
      pl_downstream_deemph_source              => '0',
      cfg_err_aer_headerlog                    => (others => '0'),
      cfg_aer_interrupt_msgnum                 => (others => '0'),
      cfg_err_aer_headerlog_set                => open,
      cfg_aer_ecrc_check_en                    => open,
      cfg_aer_ecrc_gen_en                      => open,
      cfg_vc_tcvc_map                          => open,
      config_gen_req                           => config_gen_req
   );

end architecture;



-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_pcie_mm_s_pkg.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI slave read bridge. 
--                   
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_pcie_mm_s_pkg.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;

--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------



package axi_pcie_mm_s_pkg is

   --type tag_len_array is array (0 to 7, 0 to 31) of std_logic_vector(18 downto 0);
   --type tag_len_index_array is array (0 to 7) of integer range 0 to 32;
   type cpl_addr_count_bit_array is array (0 to 7) of std_logic_vector(0 to 31);
   type tag_cpl_status_clr_array is array (0 to 7) of std_logic_vector(0 to 31);
   type first_word_offset_array is array (0 to 7) of integer range 0 to 3;
   type rresp_array is array (0 to 3) of std_logic_vector(2 downto 0);
   type slwrreqpending_array is array (0 to 3) of std_logic_vector(1 downto 0);
   type tlplength_array is array (0 to 3) of std_logic_vector(9 downto 0);
   type tlpaddrl_array is array (0 to 3) of std_logic_vector(31 downto 0);
   type barhit_array is array (0 to 3) of std_logic_vector(2 downto 0);
   type cplpendcpl_array is array (0 to 3) of std_logic;
   type wrpend_array is array (0 to 3) of std_logic_vector(3 downto 0);

   function log2(x : natural) return integer;

end package;

package body axi_pcie_mm_s_pkg is

-------------------------------------------------------------------------------
-- Function log2 -- returns number of bits needed to encode x choices
--   x = 0  returns 0
--   x = 1  returns 0
--   x = 2  returns 1
--   x = 4  returns 2, etc.
-------------------------------------------------------------------------------
--
function log2(x : natural) return integer is
   variable i  : integer := 0; 
   variable val: integer := 1;
begin 
   if x = 0 then return 0;
   else
     for j in 0 to 29 loop -- for loop for XST 
       if val >= x then null; 
       else
         i := i+1;
         val := val*2;
       end if;
     end loop;
   -- Fix per CR520627  XST was ignoring this anyway and printing a  
   -- Warning in SRP file. This will get rid of the warning and not
   -- impact simulation.  
   -- synthesis translate_off
     assert val >= x
       report "Function log2 received argument larger" &
              " than its capability of 2^30. "
       severity failure;
   -- synthesis translate_on
     return i;
   end if;  
end function log2; 
 
end package body axi_pcie_mm_s_pkg;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_mm_masterbridge_rd.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge read function
-- on the AXI memory map.
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_mm_masterbridge_rd.vhd
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

--library AMDCoreLib;
--use AMDCoreLib.all;
--library UNISIM;
--use UNISIM.VComponents.all;

entity axi_mm_masterbridge_rd is
   generic(
      --Family Generics
      C_FAMILY                : string;
      C_M_AXI_ADDR_WIDTH      : integer;
      C_M_AXI_DATA_WIDTH      : integer;
      C_PCIEBAR_NUM           : integer;
      C_PCIEBAR_AS            : integer;
      C_PCIEBAR_LEN_0         : integer;
      C_PCIEBAR2AXIBAR_0      : std_logic_vector;
      C_PCIEBAR2AXIBAR_0_SEC  : integer;
      C_PCIEBAR_LEN_1         : integer;
      C_PCIEBAR2AXIBAR_1      : std_logic_vector;
      C_PCIEBAR2AXIBAR_1_SEC  : integer;
      C_PCIEBAR_LEN_2         : integer;
      C_PCIEBAR2AXIBAR_2      : std_logic_vector;
      C_PCIEBAR2AXIBAR_2_SEC  : integer
      );
   port(
      --AXI Global
      aclk            : in  std_logic; --meaningful port name
      reset           : in  std_logic; --meaningful port name
      -- AXI Master Read Address Channel
      m_axi_araddr     : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      m_axi_arlen      : out std_logic_vector(7 downto 0); --meaningful port name
      m_axi_arsize     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_arburst    : out std_logic_vector(1 downto 0); --meaningful port name
      m_axi_arprot     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_arvalid    : out std_logic; --meaningful port name
      m_axi_arready    : in  std_logic; --meaningful port name
      m_axi_arlock     : out std_logic; --meaningful port name
      m_axi_arcache    : out std_logic_vector(3 downto 0); --meaningful port name
      -- AXI Master Read Data Channel
      m_axi_rdata      : in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axi_rresp      : in  std_logic_vector(1 downto 0); --meaningful port name
      m_axi_rlast      : in  std_logic; --meaningful port name
      m_axi_rvalid     : in  std_logic; --meaningful port name
      m_axi_rready     : out std_logic; --meaningful port name
      --Master Bridge Interrupt Strobes
      master_int      : out std_logic_vector(1 downto 0); --meaningful port name
      --Internal Interface
      rdreq           : in std_logic; --meaningful port name
      rresp           : out rresp_array; --meaningful port name
      almost_full     : in  std_logic; --meaningful port name
      dataen          : out std_logic; --meaningful port name
      tlpaddrl        : in  tlpaddrl_array; --meaningful port name
      tlplength       : in  tlplength_array; --meaningful port name
      din             : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      barhit          : in  barhit_array; --meaningful port name
      blk_lnk_up      : in  std_logic; --meaningful port name
      --Internal Interface Ordering
      slwrreqpend     : in  std_logic_vector(1 downto 0); --meaningful port name
      slwrreqpending  : out slwrreqpending_array; --meaningful port name
      compready       : out std_logic_vector(2 downto 0); --meaningful port name
      addrstreampipeline  : out std_logic_vector(2 downto 0); -- meaningful port name
      s_axi_awvalid   : in std_logic;
      rdtargetpipeline    : in  std_logic_vector(2 downto 0); --meaningful port name
      master_wr_idle      : in  std_logic --meaningful port name
      );
end axi_mm_masterbridge_rd;

architecture behavioral of axi_mm_masterbridge_rd is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

type axi_rd_master_addr_states is (idle,
                                   pcietlpinfo);

signal rdaddrsmsig         : axi_rd_master_addr_states;
type axi_rd_master_data_states is (idle,
                                   datatransfer);

signal rddatasmsig         : axi_rd_master_data_states;


signal m_axi_araddr1, m_axi_araddr2, m_axi_araddr3, m_axi_araddr4 : std_logic_vector(31 downto 0);
signal m_axi_arlen1, m_axi_arlen2, m_axi_arlen3, m_axi_arlen4     : std_logic_vector(7 downto 0);


type vector_array_type6 is array (0 to 3) of std_logic_vector(1 downto 0);
signal datatxpertlp_ram         : vector_array_type6;

type vector_array_type3 is array (0 to 3) of std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
signal m_axi_araddrtemp         : vector_array_type3;
type vector_array_type4 is array (0 to 3) of std_logic_vector(9 downto 0);
signal m_axi_arlentemp          : vector_array_type4;
type vector_array_type5 is array (0 to 3) of std_logic_vector(2 downto 0);
signal m_axi_awsizetemp         : vector_array_type5;

signal datatxpertlp             : std_logic_vector(1 downto 0);
signal rrespsig                 : std_logic_vector(1 downto 0);
signal firstdwen                : std_logic;
signal addrspipeline            : std_logic_vector(2 downto 0);
signal addrmmpipeline           : std_logic_vector(2 downto 0);
signal datammpipeline           : std_logic_vector(2 downto 0);
signal splitcnt, splitcntr      : std_logic_vector(1 downto 0);
signal m_axi_arvalid_sig        : std_logic;
signal m_axi_rdatatemp64        : std_logic_vector(31 downto 0);
signal m_axi_rdatatemp128       : std_logic_vector(95 downto 0);
signal databeat1, single_beat   : std_logic;
signal blk_lnk_up_d             : std_logic;
signal m_axi_arprottemp         : vector_array_type5;

function log2 (x : positive) return natural is 
begin
   if x = 1 then
      return 0;
   else
      return log2 (x / 2) + 1;
   end if;
end function log2;

begin

addrstreampipeline <= addrspipeline;

axi_rd_master_addr: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         rdaddrsmsig       <= idle;
         addrmmpipeline    <= "000";
         m_axi_araddr      <= (others => '0');
         m_axi_arlen       <= (others => '0');
         m_axi_arsize      <= (others => '0');
         m_axi_arprot      <= "000";
         m_axi_arvalid_sig <= '0';
         splitcnt          <= "00";
         splitcntr         <= "00";
      else
         case rdaddrsmsig is
            when idle => 
               m_axi_araddr1 <= (others => '0');
               m_axi_araddr2 <= (others => '0');
               m_axi_araddr3 <= (others => '0');
               m_axi_araddr4 <= (others => '0');
               if addrmmpipeline /= addrspipeline and master_wr_idle = '1' then
                  rdaddrsmsig     <= pcietlpinfo;
                  m_axi_araddr1 <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)));
                  splitcnt <= m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))(9 downto 8);
                  if m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))(9) = '0' then
                     if m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))(8) = '0' then
                        m_axi_arlen1 <= m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 0);
                     else
                        m_axi_arlen1 <= x"FF";
                        m_axi_arlen2 <= 
                           conv_std_logic_vector(conv_integer(m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))) - 256, 8);
                        if C_M_AXI_DATA_WIDTH = 32 then
                           m_axi_araddr2(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                             "100000000";
                        elsif C_M_AXI_DATA_WIDTH = 64 then
                           m_axi_araddr2(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                             "1000000000";
                        else
                           m_axi_araddr2(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                             "10000000000";
                        end if;
                     end if;
                  else
                     m_axi_arlen1 <= x"FF";
                     m_axi_arlen2 <= x"FF";
                     if C_M_AXI_DATA_WIDTH = 32 then
                        m_axi_araddr2(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                          "100000000";
                        m_axi_araddr3(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                          "1000000000";
                        -- coverage off
                     elsif C_M_AXI_DATA_WIDTH = 64 then
                        m_axi_araddr2(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                          "1000000000";
                        m_axi_araddr3(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                          "10000000000";
                     else
                        m_axi_araddr2(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                          "10000000000";
                        m_axi_araddr3(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                          "100000000000";
                     end if;
                        -- coverage on
                     if m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))(8) = '0' then
                        m_axi_arlen3 <= 
                           conv_std_logic_vector(conv_integer(m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))) - 512, 8);
                     else
                        m_axi_arlen3 <= x"FF";
                        m_axi_arlen4 <= 
                           conv_std_logic_vector(conv_integer(m_axi_arlentemp(conv_integer(addrmmpipeline(1 downto 0)))) - 768, 8);
                        if C_M_AXI_DATA_WIDTH = 32 then
                           m_axi_araddr4(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                             "1100000000";
                        -- coverage off
                        elsif C_M_AXI_DATA_WIDTH = 64 then
                           m_axi_araddr4(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                             "11000000000";
                        else
                           m_axi_araddr4(31 downto 2) <= m_axi_araddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(31 downto 2) + 
                             "110000000000";
                        end if;
                        -- coverage on
                     end if;
                  end if;
               else
                  rdaddrsmsig       <= idle;
                  m_axi_araddr      <= (others => '0');
                  m_axi_arlen       <= (others => '0');
                  m_axi_arsize      <= (others => '0');
                  m_axi_arprot      <= "000";
                  m_axi_arvalid_sig     <= '0';
               end if;

            when pcietlpinfo => 
               m_axi_arvalid_sig <= '1';
               if splitcntr = "00" then
                  m_axi_araddr <= m_axi_araddr1;
                  m_axi_arlen  <= m_axi_arlen1;
               elsif splitcntr = "01" then
                  m_axi_araddr <= m_axi_araddr2;
                  m_axi_arlen  <= m_axi_arlen2;
               elsif splitcntr = "10" then
                  m_axi_araddr <= m_axi_araddr3;
                  m_axi_arlen  <= m_axi_arlen3;
               else
                  m_axi_araddr <= m_axi_araddr4;
                  m_axi_arlen  <= m_axi_arlen4;
               end if;
               m_axi_arsize  <= m_axi_awsizetemp(conv_integer(addrmmpipeline(1 downto 0)));
               m_axi_arprot  <= m_axi_arprottemp(conv_integer(addrmmpipeline(1 downto 0)));
               if m_axi_arready = '1' and m_axi_arvalid_sig = '1' then
                  if splitcntr /= splitcnt then
                     rdaddrsmsig   <= pcietlpinfo;
                     splitcntr <= splitcntr + 1;
                     m_axi_arvalid_sig <= '0';
                  else
                     rdaddrsmsig   <= idle;
                     addrmmpipeline <= addrmmpipeline + 1;
                     m_axi_arvalid_sig <= '0';
                     splitcntr <= "00";
                  end if;
               end if;
               -- CR 655332
               -- Flush the request which is not received by target interface after link down event
               -- 655644
               -- Once ARVALID once asserted, will remain asserted unless until 
               -- it gets ARREADY signal
               if blk_lnk_up = '0' and m_axi_arvalid_sig = '0'  and splitcntr = "00" then
                  m_axi_arvalid_sig <= '0';
                  rdaddrsmsig       <= idle;
                  splitcntr         <= "00";
               end if;
            
            -- coverage off
            when others =>
               rdaddrsmsig <= idle;
            -- coverage on
         end case;
         --if blk_lnk_up = '0' then -- flush next read req
         --   addrmmpipeline <= addrspipeline;
         --end if;
      end if;
   end if;
end process;

data_width_32: if C_M_AXI_DATA_WIDTH = 32 generate
axi_wr_master_data: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_rready <= '0';
         rddatasmsig     <= idle;
         datammpipeline  <= (others => '0');
         rrespsig <= (others => '0');
         din <= (others => '0');
         dataen <= '0';
         datatxpertlp     <= (others => '0');
         master_int <= "00";
         single_beat <= '0';
      else
         case rddatasmsig is
            when idle =>
               m_axi_rready <= '0';
               dataen <= '0';
               master_int <= "00";
               if datammpipeline /= addrspipeline or datammpipeline(1 downto 0) /= rdtargetpipeline(1 downto 0) then
                  rresp(conv_integer(datammpipeline(1 downto 0))) <= (others => '0');
               end if;
               if datammpipeline /= addrspipeline then
                  rddatasmsig   <= datatransfer;
                  datatxpertlp <= datatxpertlp_ram(conv_integer(datammpipeline(1 downto 0)));
                  rrespsig <= (others => '0');
                  dataen <= '1';
                  single_beat <= '1';
               else
                  rddatasmsig <= idle;
                  dataen <= '0';
               end if;
            
            when datatransfer  =>
               single_beat <= '0';
               m_axi_rready <= not(almost_full);
               if almost_full = '0' then
                  if m_axi_rvalid = '1' then
                     din <= m_axi_rdata;
                     rrespsig(0) <= m_axi_rresp(0) or rrespsig(0);
                     rrespsig(1) <= m_axi_rresp(1) or rrespsig(1);
                     if m_axi_rlast = '1' then
                        if datatxpertlp /= "00" then
                           datatxpertlp <= datatxpertlp - 1;
                           rddatasmsig   <= datatransfer;
                        else
                           rddatasmsig <= idle;
                           m_axi_rready <= single_beat;
                           dataen <= single_beat;
                           datammpipeline <= datammpipeline + 1;
                           rresp(conv_integer(datammpipeline(1 downto 0))) <= 
                              '1' & (m_axi_rresp(1) or rrespsig(1)) & (m_axi_rresp(0) or rrespsig(0));
                           master_int(1) <= (m_axi_rresp(1) or rrespsig(1)) and not(m_axi_rresp(0) or rrespsig(0));
                           master_int(0) <= (m_axi_rresp(1) or rrespsig(1)) and (m_axi_rresp(0) or rrespsig(0));
                           slwrreqpending(conv_integer(datammpipeline(1 downto 0))) <= slwrreqpend + conv_integer(s_axi_awvalid);
                        end if;
                     end if;
                  end if;
               end if;
            
            -- coverage off
            when others =>
               rddatasmsig <= idle;
            -- coverage on
         end case;
         if blk_lnk_up = '0' then
           rresp <= (others => (others => '0'));
         end if;
      end if;
   end if;
end process;
end generate;

data_width_64: if C_M_AXI_DATA_WIDTH = 64 generate
axi_wr_master_data: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_rready <= '0';
         rddatasmsig     <= idle;
         datammpipeline  <= (others => '0');
         rrespsig <= (others => '0');
         m_axi_rdatatemp64 <= (others => '0');
         databeat1 <= '0';
         din <= (others => '0');
         dataen <= '0';
         datatxpertlp <= (others => '0');
         master_int <= "00";
         single_beat <= '0';
      else
         case rddatasmsig is
            when idle =>
               m_axi_rready <= '0';
               dataen <= '0';
               master_int <= "00";
               if datammpipeline /= addrspipeline or datammpipeline(1 downto 0) /= rdtargetpipeline(1 downto 0) then
                  rresp(conv_integer(datammpipeline(1 downto 0))) <= (others => '0');
               end if;
               if datammpipeline /= addrspipeline then
                  rddatasmsig   <= datatransfer;
                  datatxpertlp <= datatxpertlp_ram(conv_integer(datammpipeline(1 downto 0)));
                  rrespsig <= (others => '0');
                  dataen <= '1';
                  databeat1 <= '1';
                  single_beat <= '1';
               else
                  rddatasmsig <= idle;
                  dataen <= '0';
               end if;
            
            when datatransfer  =>
               single_beat <= '0';
               m_axi_rready <= not(almost_full);
               if almost_full = '0' then
                  if m_axi_rvalid = '1' then
                     din <= m_axi_rdata;
                     rrespsig(0) <= m_axi_rresp(0) or rrespsig(0);
                     rrespsig(1) <= m_axi_rresp(1) or rrespsig(1);
                     if m_axi_rlast = '1' then
                        if datatxpertlp /= "00" then
                           datatxpertlp <= datatxpertlp - 1;
                           rddatasmsig   <= datatransfer;
                        else
                           rddatasmsig <= idle;
                           m_axi_rready <= single_beat;
                           dataen <= single_beat;
                           datammpipeline <= datammpipeline + 1;
                           rresp(conv_integer(datammpipeline(1 downto 0))) <= 
                              '1' & (m_axi_rresp(1) or rrespsig(1)) & (m_axi_rresp(0) or rrespsig(0));
                           master_int(1) <= (m_axi_rresp(1) or rrespsig(1)) and not(m_axi_rresp(0) or rrespsig(0));
                           master_int(0) <= (m_axi_rresp(1) or rrespsig(1)) and (m_axi_rresp(0) or rrespsig(0));
                           slwrreqpending(conv_integer(datammpipeline(1 downto 0))) <= slwrreqpend + conv_integer(s_axi_awvalid);
                        end if;
                     end if;
                  end if;
               end if;
            
            -- coverage off
            when others =>
               rddatasmsig <= idle;
            -- coverage on
         end case;
         if blk_lnk_up = '0' then
           rresp <= (others => (others => '0'));
         end if;
      end if;
   end if;
end process;
end generate;

data_width_128: if C_M_AXI_DATA_WIDTH = 128 generate
axi_wr_master_data: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_rready <= '0';
         rddatasmsig     <= idle;
         datammpipeline  <= (others => '0');
         rrespsig <= (others => '0');
         m_axi_rdatatemp128 <= (others => '0');
         databeat1 <= '0';
         din <= (others => '0');
         dataen <= '0';
         datatxpertlp <= (others => '0');
         master_int <= "00";
         single_beat <= '0';
      else
         case rddatasmsig is
            when idle =>
               m_axi_rready <= '0';
               dataen <= '0';
               master_int <= "00";
               if datammpipeline /= addrspipeline or datammpipeline(1 downto 0) /= rdtargetpipeline(1 downto 0) then
                  rresp(conv_integer(datammpipeline(1 downto 0))) <= (others => '0');
               end if;
               if datammpipeline /= addrspipeline then
                  rddatasmsig   <= datatransfer;
                  datatxpertlp <= datatxpertlp_ram(conv_integer(datammpipeline(1 downto 0)));
                  rrespsig <= (others => '0');
                  dataen <= '1';
                  databeat1 <= '1';
                  single_beat <= '1';
               else
                  rddatasmsig <= idle;
                  dataen <= '0';
               end if;
            
            when datatransfer  =>
               single_beat <= '0';
               m_axi_rready <= not(almost_full);
               if almost_full = '0' then
                  if m_axi_rvalid = '1' then
                     din <= m_axi_rdata;
                     rrespsig(0) <= m_axi_rresp(0) or rrespsig(0);
                     rrespsig(1) <= m_axi_rresp(1) or rrespsig(1);
                     if m_axi_rlast = '1' then
                        if datatxpertlp /= "00" then
                           datatxpertlp <= datatxpertlp - 1;
                           rddatasmsig   <= datatransfer;
                        else
                           rddatasmsig <= idle;
                           m_axi_rready <= single_beat;
                           dataen <= single_beat;
                           datammpipeline <= datammpipeline + 1;
                           rresp(conv_integer(datammpipeline(1 downto 0))) <= 
                              '1' & (m_axi_rresp(1) or rrespsig(1)) & (m_axi_rresp(0) or rrespsig(0));
                           master_int(1) <= (m_axi_rresp(1) or rrespsig(1)) and not(m_axi_rresp(0) or rrespsig(0));
                           master_int(0) <= (m_axi_rresp(1) or rrespsig(1)) and (m_axi_rresp(0) or rrespsig(0));
                           slwrreqpending(conv_integer(datammpipeline(1 downto 0))) <= slwrreqpend + conv_integer(s_axi_awvalid);
                        end if;
                     end if;
                  end if;
               end if;
            
            -- coverage off
            when others =>
               rddatasmsig <= idle;
            -- coverage on
         end case;
         if blk_lnk_up = '0' then
           rresp <= (others => (others => '0'));
         end if;
      end if;
   end if;
end process;
end generate;

AddrTranslation: process(aclk)
   variable AddrVar : std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
   variable ARProtVar : std_logic_vector(2 downto 0);
begin
   if rising_edge(aclk) then
      if reset = '0' then
         AddrVar           := (others => '0');
         addrspipeline     <= "000";
         blk_lnk_up_d      <= '0';
      else
         if rdreq = '1' then
            for i in 0 to C_PCIEBAR_NUM-1 loop
               if barhit(conv_integer(addrspipeline(1 downto 0)))(i) = '1' then 
                  --if i < C_PCIEBAR_NUM then
                     if i = 0 then
                        AddrVar := C_PCIEBAR2AXIBAR_0(0 to C_M_AXI_ADDR_WIDTH-C_PCIEBAR_LEN_0-1) & 
                           tlpaddrl(conv_integer(addrspipeline(1 downto 0)))(C_PCIEBAR_LEN_0-1 downto 0);
                        if C_PCIEBAR2AXIBAR_0_SEC = 1 then
                           ARProtVar := "000"; -- "normal secure data" accesses only
                        else
                           ARProtVar := "010"; -- "normal non-secure data" accesses only
                        end if;
                     end if;
                     if i = 1 then
                        AddrVar := C_PCIEBAR2AXIBAR_1(0 to C_M_AXI_ADDR_WIDTH-C_PCIEBAR_LEN_1-1) & 
                           tlpaddrl(conv_integer(addrspipeline(1 downto 0)))(C_PCIEBAR_LEN_1-1 downto 0);
                        if C_PCIEBAR2AXIBAR_1_SEC = 1 then
                           ARProtVar := "000"; -- "normal secure data" accesses only
                        else
                           ARProtVar := "010"; -- "normal non-secure data" accesses only
                        end if;
                     end if;
                     if i = 2 then
                        AddrVar := C_PCIEBAR2AXIBAR_2(0 to C_M_AXI_ADDR_WIDTH-C_PCIEBAR_LEN_2-1) & 
                           tlpaddrl(conv_integer(addrspipeline(1 downto 0)))(C_PCIEBAR_LEN_2-1 downto 0);
                        if C_PCIEBAR2AXIBAR_2_SEC = 1 then
                           ARProtVar := "000"; -- "normal secure data" accesses only
                        else
                           ARProtVar := "010"; -- "normal non-secure data" accesses only
                        end if;
                     end if;
                  --end if;
               end if;
            end loop;
               m_axi_araddrtemp(conv_integer(addrspipeline(1 downto 0))) <= AddrVar;
               m_axi_arprottemp(conv_integer(addrspipeline(1 downto 0)))  <= ARProtVar;
               if tlplength(conv_integer(addrspipeline(1 downto 0))) /= "0000000001" then 
                 --workaround for 1DW requests when bus width set to 64
                  m_axi_awsizetemp(conv_integer(addrspipeline(1 downto 0))) <= conv_std_logic_vector(Log2(C_M_AXI_DATA_WIDTH/8),3);
               else
                  m_axi_awsizetemp(conv_integer(addrspipeline(1 downto 0))) <= "010";
               end if;
               if C_M_AXI_DATA_WIDTH = 32 then
                  m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <=  tlplength(conv_integer(addrspipeline(1 downto 0)))-1;
                  datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                     conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1), 10)(9 downto 8);
               else
                  if C_M_AXI_DATA_WIDTH = 64 then
                     if conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1) mod 2 = 1 and AddrVar(2) = '1' then
                        m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                           conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/2 + 1, 10);
                        datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                          conv_std_logic_vector(conv_integer(tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/2 + 
                            1, 10)(9 downto 8);
                     else
                        m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                           conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/2, 10);
                        datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                           conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/2, 
                             10)(9 downto 8);
                     end if;
                  else
                     case (conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1) mod 4) is
                     when 3 =>
                        if AddrVar(3 downto 2) = "00" then
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 
                                10)(9 downto 8);
                        else
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4 + 
                                1, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4 + 
                                1, 10)(9 downto 8);
                        end if;
                     when 0 =>
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 
                                10)(9 downto 8);
                     when 1 =>
                        if AddrVar(3 downto 2) = "11" then
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4 + 1, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4 + 
                                1, 10)(9 downto 8);
                        else
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 
                                10)(9 downto 8);
                        end if;
                     when 2 =>
                        if AddrVar(3) = '1' then
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4 + 1, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4 + 
                                1, 10)(9 downto 8);
                        else
                           m_axi_arlentemp(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 10);
                           datatxpertlp_ram(conv_integer(addrspipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer( tlplength(conv_integer(addrspipeline(1 downto 0)))-1)/4, 
                                10)(9 downto 8);
                        end if;
                     -- coverage off
                     when others =>
                     -- coverage on
                     end case;
                  end if;
               end if;
               addrspipeline <= addrspipeline + 1;

         end if;
         blk_lnk_up_d <= blk_lnk_up;
         if blk_lnk_up_d = '1' and blk_lnk_up = '0' then -- flush next read req
           -- CR 655332
           -- Just before link down transition, if any pending read request is accepted by target interface
           -- then we should expect data for the same to flush out
            if m_axi_arvalid_sig = '1' or (m_axi_arvalid_sig = '0' and splitcntr /= "00") then
               addrspipeline <= addrmmpipeline + 1;
            else
               addrspipeline <= addrmmpipeline;
            end if;
         end if;
      end if;
   end if;
end process;


m_axi_arburst <= "01"; --INCR only
m_axi_arcache <= "0011"; --cacheable & bufferable, but do not allocate
m_axi_arlock  <= '0';

m_axi_arvalid <= m_axi_arvalid_sig;
compready <= datammpipeline;

end behavioral;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_mm_masterbridge_wr.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge write function
-- on the AXI memory map.
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_mm_masterbridge_wr.vhd
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity axi_mm_masterbridge_wr is
   generic(
      --Family Generics
      C_FAMILY                : string;
      C_M_AXI_ADDR_WIDTH      : integer;
      C_M_AXI_DATA_WIDTH      : integer;
      C_PCIEBAR_NUM           : integer;
      C_PCIEBAR_AS            : integer;
      C_PCIEBAR_LEN_0         : integer;
      C_PCIEBAR2AXIBAR_0      : std_logic_vector;
      C_PCIEBAR2AXIBAR_0_SEC  : integer;
      C_PCIEBAR_LEN_1         : integer;
      C_PCIEBAR2AXIBAR_1      : std_logic_vector;
      C_PCIEBAR2AXIBAR_1_SEC  : integer;
      C_PCIEBAR_LEN_2         : integer;
      C_PCIEBAR2AXIBAR_2      : std_logic_vector;
      C_PCIEBAR2AXIBAR_2_SEC  : integer
      );
   port(
      --AXI Global
      aclk            : in  std_logic; --meaningful port name
      reset           : in  std_logic; --meaningful port name
      --AXI master Write Address Channel
      m_axi_awaddr    : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      m_axi_awlen     : out std_logic_vector(7 downto 0); --meaningful port name
      m_axi_awsize    : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_awburst   : out std_logic_vector(1 downto 0); --meaningful port name
      m_axi_awprot    : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_awvalid   : out std_logic; --meaningful port name
      m_axi_awready   : in std_logic; --meaningful port name
      m_axi_awlock    : out std_logic; --meaningful port name
      m_axi_awcache   : out std_logic_vector(3 downto 0); --meaningful port name
      --AXI master Write Data Channel
      m_axi_wdata     : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axi_wstrb     : out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0); --meaningful port name
      m_axi_wlast     : out std_logic; --meaningful port name
      m_axi_wvalid    : out std_logic; --meaningful port name
      m_axi_wready    : in  std_logic; --meaningful port name
      --AXI master Write Response Channel
      m_axi_bresp     : in  std_logic_vector(1 downto 0); --meaningful port name
      m_axi_bvalid    : in  std_logic; --meaningful port name
      m_axi_bready    : out std_logic; --meaningful port name
      --Master Bridge Interrupt Strobes
      master_int      : out std_logic_vector(1 downto 0); --meaningful port name
      --Internal Interface
      wrreqset        : in  std_logic; --meaningful port name
      datacompcheck   : out std_logic; --meaningful port name (used for self testing)
      tlplength       : in  std_logic_vector(9 downto 0); --meaningful port name
      firstdwbe       : in  std_logic_vector(3 downto 0); --meaningful port name
      lastdwbe        : in  std_logic_vector(3 downto 0); --meaningful port name
      tlpaddrl        : in  std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      tlpaddrh        : in  std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name (not used)
      dout            : in  std_logic_vector(C_M_AXI_DATA_WIDTH downto 0); --meaningful port name
      rd_en           : out std_logic; --meaningful port name
      empty           : in  std_logic; --meaningful port name
      tlppipeline     : out std_logic_vector(2 downto 0); --meaningful port name
      barhit          : in  std_logic_vector(C_PCIEBAR_NUM-1 downto 0); --meaningful port name
      --Internal Interface Ordering
      wrreqcomp       : out std_logic_vector(2 downto 0) --meaningful port name
      );
end axi_mm_masterbridge_wr;

architecture behavioral of axi_mm_masterbridge_wr is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

type axi_wr_master_addr_states is (idle,
                                   pcietlpinfo);

signal wraddrsmsig         : axi_wr_master_addr_states;
type axi_wr_master_data_states is (idle,
                                   datatransfer32,
                                   datatransfer64,
                                   datatransfer128);

signal wrdatasmsig         : axi_wr_master_data_states;
type axi_wr_master_resp_states is (idle,
                                   respreport);

signal wrrespsmsig         : axi_wr_master_resp_states;


type vector_array_type4 is array (0 to 3) of std_logic_vector(1 downto 0);
signal m_axi_awaddrsttemp  : vector_array_type4;

type vector_array_type8 is array (0 to 3) of std_logic_vector(7 downto 0);
signal m_axi_awlensttemp     : vector_array_type8;

type vector_array_type7 is array (0 to 3) of std_logic_vector(3 downto 0);
signal firstdwbetemp, lastdwbetemp       : vector_array_type7;

type vector_array_type3 is array (0 to 3) of std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
signal m_axi_awaddrtemp    : vector_array_type3;
type vector_array_type5 is array (0 to 3) of std_logic_vector(7 downto 0);
signal m_axi_awlentemp     : vector_array_type5;
type vector_array_type6 is array (0 to 3) of std_logic_vector(2 downto 0);
signal m_axi_awsizetemp    : vector_array_type6;
signal firstdwen           : std_logic;
signal wrreqsetcnt     : std_logic_vector(2 downto 0);
signal tlplength_reg       : std_logic_vector(7 downto 0);
signal m_axi_awvalidsig    : std_logic;
signal m_axi_wvalidsig     : std_logic;
signal m_axi_breadysig     : std_logic;
signal addrspipeline       : std_logic_vector(2 downto 0);
signal addrmmpipeline      : std_logic_vector(2 downto 0);
signal datammpipeline      : std_logic_vector(2 downto 0);
signal respmmpipeline      : std_logic_vector(2 downto 0);
signal m_axi_awprottemp    : vector_array_type6;

function log2 (x : positive) return natural is 
begin
   if x = 1 then
      return 0;
   else
      return log2 (x / 2) + 1;
   end if;
end function log2;

begin

axi_wr_master_addr: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_awaddr      <= (others => '0');
         m_axi_awlen       <= (others => '0');
         m_axi_awsize      <= (others => '0');
         m_axi_awprot      <= "000";
         m_axi_awvalidsig  <= '0';
         wraddrsmsig       <= idle;
         addrmmpipeline    <= "000";
      else
         case wraddrsmsig is
            when idle => 
               m_axi_awvalidsig     <= '0';
               if addrmmpipeline /= addrspipeline then
                  wraddrsmsig     <= pcietlpinfo;
               else
                  m_axi_awaddr      <= (others => '0');
                  m_axi_awlen       <= (others => '0');
                  m_axi_awsize      <= (others => '0');
                  m_axi_awprot      <= "000";
               end if;

            when pcietlpinfo => 
               m_axi_awvalidsig <= '1';
               m_axi_awaddr  <= m_axi_awaddrtemp(conv_integer(addrmmpipeline(1 downto 0)));
               if C_M_AXI_DATA_WIDTH = 32 then
                  m_axi_awlen   <= m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)));
               elsif C_M_AXI_DATA_WIDTH = 64 then
                  if m_axi_awaddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(2) = '1' and 
                     m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(0) = '1' then
                     m_axi_awlen   <= 
                        '0' & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 1) + 
                           "00000001";
                  else
                     m_axi_awlen   <= 
                        '0' & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 1);
                  end if;
               else
                  case (m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(1 downto 0)) is
                  when "11" =>
                     if m_axi_awaddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(3 downto 2) = "00" then
                        m_axi_awlen   <= 
                           "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2);
                     else
                        m_axi_awlen   <= 
                           "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2) + 
                              "00000001";
                     end if;
                  when "00" =>
                     m_axi_awlen   <= 
                        "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2);
                  when "01" =>
                     if m_axi_awaddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(3 downto 2) = "11" then
                        m_axi_awlen   <= 
                           "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2) + 
                              "00000001";
                     else
                        m_axi_awlen   <= 
                           "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2);
                     end if;
                  when "10" =>
                     if m_axi_awaddrtemp(conv_integer(addrmmpipeline(1 downto 0)))(3) = '1' then
                        m_axi_awlen   <= 
                           "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2) + 
                              "00000001";
                     else
                        m_axi_awlen   <= 
                           "00" & m_axi_awlentemp(conv_integer(addrmmpipeline(1 downto 0)))(7 downto 2);
                     end if;
                  when others =>
                  end case;
               end if;
               m_axi_awsize  <= m_axi_awsizetemp(conv_integer(addrmmpipeline(1 downto 0)));
               m_axi_awprot  <= m_axi_awprottemp(conv_integer(addrmmpipeline(1 downto 0)));
               if m_axi_awready = '1' and m_axi_awvalidsig = '1' then
                  wraddrsmsig   <= idle;
                  addrmmpipeline <= addrmmpipeline + 1;
                  m_axi_awvalidsig <= '0';
               end if;

            -- coverage off
            when others => 
               wraddrsmsig <= idle;
            -- coverage on
         end case;
      end if;
   end if;
end process;

data_width_32: if C_M_AXI_DATA_WIDTH = 32 generate
axi_wr_master_data: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_wvalidsig <= '0';
         datacompcheck   <= '0';
         tlplength_reg   <= (others => '0');
         wrdatasmsig     <= idle;
         firstdwen       <= '0';
         datammpipeline  <= (others => '0');
         m_axi_wstrb     <= (others => '0');
      else
            case wrdatasmsig is
               when idle =>
                  datacompcheck   <= '0';
                  if datammpipeline /= addrspipeline then
                     wrdatasmsig   <= datatransfer32;
                     firstdwen     <= '1';
                     m_axi_wstrb     <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                     tlplength_reg   <= m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)));
                  else
                     tlplength_reg   <= (others => '0');
                  end if;
               
               when datatransfer32  =>
                  m_axi_wvalidsig <= not(empty);
                  if empty = '0' then
                     if m_axi_wready = '1' then
                        if  m_axi_wvalidsig = '1' then
                           if firstdwen = '1' then
                              firstdwen   <= '0';
                           end if;
                           if dout(C_M_AXI_DATA_WIDTH) = '1' then
                              wrdatasmsig <= idle;
                              m_axi_wvalidsig <= '0';
                              datacompcheck <= '1';
                              datammpipeline <= datammpipeline + 1;
                           end if;
                           if tlplength_reg = x"01" then
                              m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                           else
                              m_axi_wstrb     <= (others => '1');
                           end if;
                           tlplength_reg <= tlplength_reg - 1;
                        end if;
                     end if;
                  end if;
               
               -- coverage off
               when others =>
                  wrdatasmsig <= idle;
               -- coverage on
            end case;
      end if;
   end if;
end process;
end generate;
         
data_width_64: if C_M_AXI_DATA_WIDTH = 64 generate
axi_wr_master_data: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_wvalidsig <= '0';
         datacompcheck   <= '0';
         tlplength_reg   <= (others => '0');
         wrdatasmsig     <= idle;
         firstdwen       <= '0';
         datammpipeline  <= (others => '0');
         m_axi_wstrb     <= (others => '0');
      else
            case wrdatasmsig is
               when idle            => 
                  datacompcheck   <= '0';
                  if datammpipeline /= addrspipeline then
                     wrdatasmsig   <= datatransfer64;
                     firstdwen     <= '1';
                     if m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0))) = "00000000" then
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" or 
                           m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= x"0" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        end if;
                     elsif m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0))) = "00000001" then
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" or 
                           m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        end if;
                     else
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" or 
                           m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= x"F" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        end if;
                     end if;
                     if (m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" or 
                        m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "11") and 
                           m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(0) = '1' then
                        tlplength_reg   <= 
                           '0' & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 1) + 
                              "00000001";
                     else
                        tlplength_reg   <= 
                           '0' & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 1);
                     end if;
                  else
                     tlplength_reg   <= (others => '0');
                  end if;
               
               when datatransfer64  => 
                  m_axi_wvalidsig <= not(empty);
                  if empty = '0' then
                     if m_axi_wready = '1' then
                        if  m_axi_wvalidsig = '1' then
                           if firstdwen = '1' then
                              firstdwen   <= '0';
                           end if;
                           if dout(C_M_AXI_DATA_WIDTH) = '1' then
                              wrdatasmsig <= idle;
                              m_axi_wvalidsig <= '0';
                              datacompcheck <= '1';
                              datammpipeline <= datammpipeline + 1;
                           end if;
                           if tlplength_reg = x"01" then
                              if m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(0) = '1' then
                                 if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" or 
                                    m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                                    m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F";
                                 else
                                    m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                                 end if;
                              else
                                 if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" or 
                                    m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                                    m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                                 else
                                    m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F";
                                 end if;
                              end if;
                           else
                              m_axi_wstrb <= (others => '1');
                           end if;
                           tlplength_reg <= tlplength_reg - 1;
                        end if;
                     end if;
                  end if;

               -- coverage off
               when others =>
                  wrdatasmsig <= idle;
               -- coverage on
            end case;
      end if;
   end if;
end process;
end generate;
         
data_width_128: if C_M_AXI_DATA_WIDTH = 128 generate
axi_wr_master_data: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_wvalidsig <= '0';
         datacompcheck   <= '0';
         tlplength_reg   <= (others => '0');
         wrdatasmsig     <= idle;
         firstdwen       <= '0';
         datammpipeline  <= (others => '0');
         m_axi_wstrb     <= (others => '0');
      else
            case wrdatasmsig is
               when idle            => 
                  datacompcheck   <= '0';
                  if datammpipeline /= addrspipeline then
                     wrdatasmsig   <= datatransfer128;
                     firstdwen     <= '1';
                     case (conv_integer(m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0))))) is
                     when 0 =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                           m_axi_wstrb <= x"000" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                           m_axi_wstrb <= x"00" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= x"0" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"00";
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"000";
                        end if;
                     when 1 =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                           m_axi_wstrb <= x"00" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                           m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"00";
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"000";
                        end if;
                     when 2 =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                           m_axi_wstrb <= x"0"& lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F" & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                           m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F" & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= x"F" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"00";
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"000";
                        end if;
                     when 3 =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                           m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FF" & 
                              firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                           m_axi_wstrb <= x"FF" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= x"F" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"00";
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"000";
                        end if;
                     when others =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                           m_axi_wstrb <= x"FFF" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                           m_axi_wstrb <= x"FF" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"0";
                        elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                           m_axi_wstrb <= x"F" & firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"00";
                        else
                           m_axi_wstrb <= firstdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"000";
                        end if;
                     end case;
                     case (m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(1 downto 0)) is
                     when "11" =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                           tlplength_reg   <= 
                              "00" & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 2);
                        else
                           tlplength_reg   <= 
                              "00" & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 2)
                                 + "00000001";
                        end if;
                     when "00" =>
                        tlplength_reg   <= 
                           "00" & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 2);
                     when "01" =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "11" then
                           tlplength_reg   <= 
                              "00" & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 2)
                                 + "00000001";
                        else
                           tlplength_reg   <= 
                              conv_std_logic_vector(conv_integer(m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0))))/4, 8);
                        end if;
                     when "10" =>
                        if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" or 
                           m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "11" then
                           tlplength_reg   <= 
                              "00" & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 2)
                                 + "00000001";
                        else
                           tlplength_reg <= 
                              "00" & m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(7 downto 2);
                        end if;
                     -- coverage off
                     when others =>
                     -- coverage on
                     end case;
                  else
                     tlplength_reg   <= (others => '0');
                  end if;
               
               when datatransfer128 => 
                  m_axi_wvalidsig <= not(empty);
                  if empty = '0' then
                     if m_axi_wready = '1' then
                        if  m_axi_wvalidsig = '1' then
                           if firstdwen = '1' then
                              firstdwen   <= '0';
                           end if;
                           if dout(C_M_AXI_DATA_WIDTH) = '1' then
                              wrdatasmsig <= idle;
                              m_axi_wvalidsig <= '0';
                              datacompcheck <= '1';
                              datammpipeline <= datammpipeline + 1;
                           end if;
                           if tlplength_reg = x"01" then
                              case (m_axi_awlensttemp(conv_integer(datammpipeline(1 downto 0)))(1 downto 0)) is
                              when "11" =>
                                 if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                                    m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FFF";
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                                    m_axi_wstrb <= x"000" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                                    m_axi_wstrb <= x"00" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F";
                                 else
                                    m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FF";
                                 end if;
                              when "00" =>
                                 if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                                    m_axi_wstrb <= x"000" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                                    m_axi_wstrb <= x"00" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F";
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                                    m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FF";
                                 else
                                    m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FFF";
                                 end if;
                              when "01" =>
                                 if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                                    m_axi_wstrb <= x"00" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F";
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                                    m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FF";
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                                    m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FFF";
                                 else
                                    m_axi_wstrb <= x"000" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                                 end if;
                              when "10" =>
                                 if m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "00" then
                                    m_axi_wstrb <= x"0" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FF";
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "01" then
                                    m_axi_wstrb <= lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"FFF";
                                 elsif m_axi_awaddrsttemp(conv_integer(datammpipeline(1 downto 0))) = "10" then
                                    m_axi_wstrb <= x"000" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0)));
                                 else
                                    m_axi_wstrb <= x"00" & lastdwbetemp(conv_integer(datammpipeline(1 downto 0))) & x"F";
                                 end if;
                              -- coverage off
                              when others =>
                              -- coverage on
                              end case;
                           else
                              m_axi_wstrb <= (others => '1');
                           end if;
                           tlplength_reg <= tlplength_reg - 1;
                        end if;
                     end if;
                  end if;

               -- coverage off
               when others=>
                  wrdatasmsig <= idle;
               -- coverage on
            end case;
      end if;
   end if;
end process;
end generate;

axi_wr_master_resp: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         m_axi_breadysig    <= '0';
         master_int      <= "00";
         wrrespsmsig     <= idle;
         respmmpipeline  <= "000";
      else
         case wrrespsmsig is
            when idle       => 
               master_int <= "00";
               if respmmpipeline /= addrspipeline then
                  m_axi_breadysig <= '1';
                  wrrespsmsig <= respreport;
               else
                  m_axi_breadysig <= '0';
               end if;
            
            when respreport => 
               if m_axi_bvalid = '1' then
                  wrrespsmsig <= idle;
                  m_axi_breadysig <= '0';
                  if m_axi_bresp = "11" then            --DECERR
                     master_int(0) <= '1';              --Master DECERR Interrupt Strobe
                  elsif m_axi_bresp = "10" then         --SLVERR
                     master_int(1) <= '1';              --Master SLVERR Interrupt Strobe
                  end if;
                  respmmpipeline <= respmmpipeline + 1;
               end if;
            
            -- coverage off
            when others => 
               wrrespsmsig <= idle;
            -- coverage on
         end case;
      end if;
   end if;
end process;

AddrTranslation: process(aclk)
   variable AddrVar : std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
   variable AWProtVar : std_logic_vector(2 downto 0);
begin
   if rising_edge(aclk) then
      if reset = '0' then
         AddrVar           := (others => '0');
         addrspipeline     <= "000";
         AWProtVar         := (others => '0');
      else
         if wrreqset = '1' then
            for i in 0 to C_PCIEBAR_NUM-1 loop
               if barhit(i) = '1' then 
                  if i < C_PCIEBAR_NUM then
                     if i = 0 then
                        AddrVar := C_PCIEBAR2AXIBAR_0(0 to C_M_AXI_ADDR_WIDTH-C_PCIEBAR_LEN_0-1) & 
                           tlpaddrl(C_PCIEBAR_LEN_0-1 downto 0);
                        if C_PCIEBAR2AXIBAR_0_SEC = 1 then
                           AWProtVar := "000"; -- "normal secure data" accesses only
                        else
                           AWProtVar := "010"; -- "normal non-secure data" accesses only
                        end if;
                     end if;
                     if i = 1 then
                        AddrVar := C_PCIEBAR2AXIBAR_1(0 to C_M_AXI_ADDR_WIDTH-C_PCIEBAR_LEN_1-1) & 
                           tlpaddrl(C_PCIEBAR_LEN_1-1 downto 0);
                        if C_PCIEBAR2AXIBAR_1_SEC = 1 then
                           AWProtVar := "000"; -- "normal secure data" accesses only
                        else
                           AWProtVar := "010"; -- "normal non-secure data" accesses only
                        end if;
                     end if;
                     if i = 2 then
                        AddrVar := C_PCIEBAR2AXIBAR_2(0 to C_M_AXI_ADDR_WIDTH-C_PCIEBAR_LEN_2-1) & 
                           tlpaddrl(C_PCIEBAR_LEN_2-1 downto 0);
                        if C_PCIEBAR2AXIBAR_2_SEC = 1 then
                           AWProtVar := "000"; -- "normal secure data" accesses only
                        else
                           AWProtVar := "010"; -- "normal non-secure data" accesses only
                        end if;
                     end if;
                  end if;
               end if;
            end loop;
               m_axi_awaddrtemp(conv_integer(addrspipeline(1 downto 0)))               <= AddrVar;
               m_axi_awaddrsttemp(conv_integer(addrspipeline(1 downto 0))) <= AddrVar(3 downto 2);
               --if tlplength(8) = '0' then --Xilinx core would only support max payload of 256bytes for v6/s6
                  m_axi_awlentemp(conv_integer(addrspipeline(1 downto 0)))   <= tlplength(7 downto 0) - 1;
                  m_axi_awlensttemp(conv_integer(addrspipeline(1 downto 0)))   <= tlplength(7 downto 0) - 1;
               --else
               --   m_axi_awlentemp(conv_integer(addrspipeline(1 downto 0)))   <= (others => '1');
               --   m_axi_awlensttemp(conv_integer(addrspipeline(1 downto 0)))   <= (others => '1');
               --end if;
               if tlplength /= "0000000001" then --workaround for 1DW requests when bus width set to 64
                  m_axi_awsizetemp(conv_integer(addrspipeline(1 downto 0)))  <= conv_std_logic_vector(Log2(C_M_AXI_DATA_WIDTH/8),3);
               else
                  m_axi_awsizetemp(conv_integer(addrspipeline(1 downto 0))) <= "010";
               end if;
               firstdwbetemp(conv_integer(addrspipeline(1 downto 0)))     <= firstdwbe;
               lastdwbetemp(conv_integer(addrspipeline(1 downto 0)))      <= lastdwbe;
               m_axi_awprottemp(conv_integer(addrspipeline(1 downto 0)))  <= AWProtVar;
               addrspipeline <= addrspipeline + 1;
         end if;
      end if;
   end if;
end process;


Pipeline: process(aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         wrreqsetcnt <= "000";
      elsif wrreqset = '1' and m_axi_bvalid = '1' and m_axi_breadysig = '1' then
         wrreqsetcnt <= wrreqsetcnt;
      elsif wrreqset = '1' then
         wrreqsetcnt<= wrreqsetcnt + 1;
      elsif m_axi_bvalid = '1' and m_axi_breadysig = '1' then
         wrreqsetcnt<= wrreqsetcnt - 1;
      end if;
   end if;
end process;

m_axi_awvalid    <= m_axi_awvalidsig;
m_axi_bready     <= m_axi_breadysig;
m_axi_wvalid     <= 
   m_axi_wvalidsig when empty = '0' else
   '0';
tlppipeline  <= wrreqsetcnt;
rd_en            <= m_axi_wready and m_axi_wvalidsig and not(empty);
m_axi_wdata      <= 
   dout(C_M_AXI_DATA_WIDTH-1 downto 0) when datammpipeline /= addrspipeline else
   (others => '0');
m_axi_wlast      <= 
   dout(C_M_AXI_DATA_WIDTH) when datammpipeline /= addrspipeline else
   '0';

m_axi_awburst <= "01"; --INCR only
m_axi_awcache <= "0011"; --cacheable & bufferable, but do not allocate
m_axi_awlock  <= '0';

wrreqcomp <= respmmpipeline;

end behavioral;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_s_masterbridge_rd.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge read function
-- on the AXI Stream.
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_s_masterbridge_rd.vhd
--
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.conv_std_logic_vector;

entity array_arith is
      port(
      din0 : in integer range 0 to 1023;
      din1 : in integer range 0 to 1023;
      dout : out std_logic_vector(9 downto 0)
      );
end array_arith;

architecture rtl of array_arith is
      attribute DONT_TOUCH : string;
      attribute DONT_TOUCH of rtl : architecture is "true";
      signal din2 : integer range 0 to 2047;
      signal din3 : integer range 0 to 511;
      signal dout_tmp : integer range 0 to 1;
begin
      din2 <= din0 + din1;
      dout_tmp <= 0 when (din2 mod 4) = 0 else 1;
      din3 <= (din0 + din1)/4;                      
      dout <= conv_std_logic_vector(din3 + dout_tmp, 10);
end rtl;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

entity axi_s_masterbridge_rd is
   generic(
      --Family Generics
      C_FAMILY            : string := "artix7";
      C_S_AXIS_DATA_WIDTH : integer := 128;
      C_S_AXIS_USER_WIDTH : integer := 22;
      C_PCIEBAR_NUM       : integer := 1;
      C_PCIEBAR_AS        : integer := 0;
      C_TRN_NP_FC         : string  := "FALSE"
      );
   port(
      --AXI Global
      aclk             : in  std_logic; --meaningful port name
      reset            : in  std_logic; --meaningful port name
      -- AXIS Read Target Channel
      s_axis_cr_tdata  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      s_axis_cr_tstrb  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      s_axis_cr_tlast  : in  std_logic; --meaningful port name
      s_axis_cr_tvalid : in  std_logic; --meaningful port name
      s_axis_cr_tready : out std_logic; --meaningful port name
      s_axis_cr_tuser  : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      -- AXIS Completion Target Channel
      m_axis_cc_tdata  : out std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axis_cc_tstrb  : out std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      m_axis_cc_tlast  : out std_logic; --meaningful port name
      m_axis_cc_tvalid : out std_logic; --meaningful port name
      m_axis_cc_tready : in  std_logic; --meaningful port name
      m_axis_cc_tuser  : out std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --AXI Streaming Block Interface
      blk_lnk_up          : in  std_logic; --meaningful port name
      blk_dcontrol        : in  std_logic_vector(15 downto 0); --meaningful port name
      blk_bus_number      : in  std_logic_vector(7 downto 0); --meaningful port name
      blk_device_number   : in  std_logic_vector(4 downto 0); --meaningful port name
      blk_function_number : in  std_logic_vector(2 downto 0); --meaningful port name
      --Internal Interface
      rresp           : in  rresp_array; --meaningful port name
      rdreq           : out std_logic; --meaningful port name
      empty           : in  std_logic; --meaningful port name
      dout            : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      tlpaddrl_out    : out tlpaddrl_array; --meaningful port name
      tlplength_out   : out tlplength_array; --meaningful port name
      rd_en           : out std_logic; --meaningful port name
      --Internal Interface Ordering
      rdtargetpipeline_out : out std_logic_vector(2 downto 0); --meaningful port name
      orrdreqpipeline : in std_logic_vector(2 downto 0); --meaningful port name
      cplpendcpl      : in  cplpendcpl_array; --meaningful port name
      wrpending       : out wrpend_array; --meaningful port name
      wrreqpend       : in  std_logic_vector(2 downto 0); --meaningful port name
      slv_write_idle  : in  std_logic; --meaningful port name
      master_wr_idle  : in  std_logic; --meaningful port name
      wrreqcomp       : in  std_logic_vector(2 downto 0); --meaningful port name
      addrstreampipeline : in std_logic_vector(2 downto 0); -- meaningful port name
      blk_lnk_up_latch_o : out std_logic; --meaningful port name
      rdndreqpipeline_o  : out std_logic_vector(2 downto 0); -- Used in NP OK mode
      rdreqpipeline_o    : out std_logic_vector(2 downto 0); -- Used in NP OK mode
      np_pkt_complete_o  : out std_logic_vector(1 downto 0); -- Used in NP Req mode. bit[1] = rdndreqpipeline; bit[0] = rdreqpipeline
      s_axis_cr_tusersig : out barhit_array --meaningful port name
      );
end axi_s_masterbridge_rd;

architecture behavioral of axi_s_masterbridge_rd is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

signal tlplength_array_val : integer range 0 to 1023;
signal rdtlpaddrl_array_val : integer range 0 to 1023;
signal rdtlpaddrltemp_array_val : integer range 0 to 1023;
signal tlplengthcntr_var_tmp : std_logic_vector(9 downto 0);
signal tlplengthcntr_tmp : std_logic_vector(9 downto 0);

type rd_master_ingress_states is (init,
                                  memrdreq,
                                  blklinkdown,
                                  throttle,
                                  throttle_nd,
                                  latch_reqid_tag_be,
                                  latchaddrh,
                                  latchaddrl);

signal rdreqsmsig                            : rd_master_ingress_states;

type cpl_master_egress_states is (idle,
                                  memcplpipeline,
                                  memcplcrtdatabeat1,
                                  blklinkdown_corruptdata,
                                  memcplcrtdatabeat2,
                                  memcpltxonedw,
                                  memcpltxdata);

signal cpltlpsmsig                           : cpl_master_egress_states;

type cplnd_master_egress_states is (idle,
                                  memcplcrtdatabeat1,
                                  memcplcrtdatabeat2,
                                  transfer_complete,
                                  memcplcrtdatabeat3);

signal cplndtlpsmsig                           : cplnd_master_egress_states;

type cpl_split_states is (idle,
                          cpldsplitcalc,
                          cpldsplitparam);

signal cpldsplitsm                           : cpl_split_states;


--byte count array (0 to 1 -> book keeping per read req, 0 to 3 -> pipeline book keeping)
type ctlpbytecount_array is array (0 to 1, 0 to 3) of std_logic_vector(11 downto 0);
signal ctlpbytecount                         : ctlpbytecount_array;

--length array (0 to 2 -> book keeping per read req, 0 to 3 -> pipeline book keeping)
-- array(0 -> ragged, 1 -> maxpayload, 3 -> residue)
type ctlplength_array is array (0 to 2, 0 to 3) of std_logic_vector(9 downto 0);
signal ctlplength                            : ctlplength_array;

type vector_array_type1 is array (0 to 3) of std_logic_vector(11 downto 0);
signal tlpbytecount, tlpndbytecount          : vector_array_type1;
signal ctlpbytecount0,ctlpbytecount1         : vector_array_type1;

type vector_array_type2 is array (0 to 3) of std_logic_vector(15 downto 0);
signal tlprequesterid, tlpcompleterid      : vector_array_type2;

type vector_array_type3 is array (0 to 3) of std_logic_vector(7 downto 0);
signal tlptag                                : vector_array_type3;

type vector_array_type4 is array (0 to 3) of std_logic_vector(6 downto 0);
signal rdtlpaddrl                            : vector_array_type4;

type vector_array_type6 is array (0 to 3) of std_logic_vector(4 downto 0);
signal cpldsplitcount                        : vector_array_type6;

type vector_array_type7 is array (0 to 3) of std_logic_vector(2 downto 0);
signal tlptc                          : vector_array_type7;

type vector_array_type9 is array (0 to 3) of std_logic_vector(1 downto 0);
signal tlpattr                       : vector_array_type9;

type vector_array_type10 is array (0 to 3) of std_logic_vector(9 downto 0);
signal tlplength                             : vector_array_type10;
signal ctlplength0, ctlplength1, ctlplength2 : vector_array_type10;

type vector_array_type11 is array (0 to 3) of std_logic_vector(31 downto 0);
signal tlpaddrl                              : vector_array_type11;

type vector_array_type12 is array (0 to 3) of std_logic_vector(15 downto 0);
signal tlpndrequesterid, tlpndcompleterid  : vector_array_type12;
type vector_array_type13 is array (0 to 3) of std_logic_vector(7 downto 0);
signal tlpndtag                              : vector_array_type13;
signal rdtlpaddrltemp                        : std_logic_vector(6 downto 0);
type vector_array_type14 is array (0 to 3) of std_logic_vector(6 downto 0);
signal rdndtlpaddrl                          : vector_array_type14;
type vector_array_type15 is array (0 to 3) of std_logic_vector(2 downto 0);
signal tlpndtc, cplndstatuscode              : vector_array_type15;
type vector_array_type16 is array (0 to 3) of std_logic_vector(1 downto 0);
signal tlpndattr                             : vector_array_type16;

signal tlpaddrlow                            : std_logic_vector(31 downto 0);
signal ctlpbytecounttemp                     : std_logic_vector(11 downto 0);
signal ctlplengthtemp                        : std_logic_vector(9 downto 0);
signal tlpbytecounttemp                      : std_logic_vector(11 downto 0);
signal tlpaddrltemp                          : std_logic_vector(31 downto 0);
signal tlpaddrhigh                           : std_logic_vector(31 downto 0);
signal requesteridsig                        : std_logic_vector(15 downto 0);
signal tagsig                                : std_logic_vector(7 downto 0);
signal cplcounter, cpldsplitcounttemp        : std_logic_vector(4 downto 0);
signal np_pkt_complete                       : std_logic_vector(1 downto 0);
signal rdreqpipeline                         : std_logic_vector(2 downto 0);
signal rdndreqpipeline                       : std_logic_vector(2 downto 0);
signal rdtargetpipeline                      : std_logic_vector(2 downto 0);
signal rdndtargetpipeline                    : std_logic_vector(2 downto 0);
signal cpltargetpipeline                     : std_logic_vector(2 downto 0);
signal cplndtargetpipeline, orcplndpipeline  : std_logic_vector(2 downto 0);
signal ctargetpipeline                       : std_logic_vector(2 downto 0);
signal rdreqpipelineincr, rdreqpipelinedecr  : std_logic;
signal rdndreqpipelineincr, rdndreqpipelinedecr  : std_logic;
signal tlptcsig                              : std_logic_vector(2 downto 0);
signal tlpepsig, tlptdsig                    : std_logic;
signal bcm, cplpacket1, firstdwen            : std_logic;
signal tlpfmtsig, tlpattrsig                 : std_logic_vector(1 downto 0);
signal tlptypesig                            : std_logic_vector(4 downto 0);
signal tlplengthsig, tlplengthcntr           : std_logic_vector(9 downto 0);
signal firstdwbesig, lastdwbesig             : std_logic_vector(3 downto 0);
signal badreadreq, zerolenreadreq            : std_logic;
signal rdndtlpaddrlow                        : std_logic_vector(6 downto 0);
signal m_axis_cc_tdatatemp64                 : std_logic_vector(31 downto 0);
signal m_axis_cc_tdatatemp128                : std_logic_vector(95 downto 0);
signal lnkdowndataflush, corruptdataflush      : std_logic;
signal blk_lnk_up_latch                        : std_logic;
signal blk_lnk_up_d                            : std_logic;
-- 2 sets of signals to send cpl's for no barhit & zero len read reqs
signal m_axis_cc_tdata_d, m_axis_cc_tdata_nd   : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
signal m_axis_cc_tstrb_d, m_axis_cc_tstrb_nd   : std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
signal m_axis_cc_tlast_d, m_axis_cc_tlast_nd   : std_logic;
signal m_axis_cc_tvalid_d, m_axis_cc_tvalid_nd : std_logic;
signal length_offset                           : std_logic_vector(11 downto 0);
signal m_axis_cc_tdata_h                       : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
signal dis_valid_d, dis_valid_nd               : std_logic;
signal data_phase, rd_en_sig, dis_rden         : std_logic;
signal wait_till_not_empty                     : std_logic;
signal s_axis_cr_tready_sig                    : std_logic;
signal totallength, linkdownflushdepth         : std_logic_vector(9 downto 0);
signal totalbytecount                          : std_logic_vector(11 downto 0);
signal s_axis_cr_tusersigtemp                  : std_logic_vector(2 downto 0);
--ordering control signals
signal rrespdelayed                            : std_logic;
signal wrpendingsig, wrpendflush               : wrpend_array;
signal cplndpendcpl                            : cplpendcpl_array;

component array_arith is
      port(
      din0 : in integer range 0 to 1023;
      din1 : in integer range 0 to 1023;
      dout : out std_logic_vector(9 downto 0)
      );
end component;


function little_to_big_endian32(datain : std_logic_vector(31 downto 0))
      return std_logic_vector is
   variable dataout : std_logic_vector(31 downto 0);
begin
   dataout := datain(7 downto 0) & datain(15 downto 8) & datain(23 downto 16) & datain(31 downto 24);
   return(dataout);
end function;

begin

ctlplength0(0)      <= ctlplength(0,0);
ctlplength0(1)      <= ctlplength(0,1);
ctlplength0(2)      <= ctlplength(0,2);
ctlplength0(3)      <= ctlplength(0,3);
ctlplength1(0)      <= ctlplength(1,0);
ctlplength1(1)      <= ctlplength(1,1);
ctlplength1(2)      <= ctlplength(1,2);
ctlplength1(3)      <= ctlplength(1,3);
ctlplength2(0)      <= ctlplength(2,0);
ctlplength2(1)      <= ctlplength(2,1);
ctlplength2(2)      <= ctlplength(2,2);
ctlplength2(3)      <= ctlplength(2,3);
ctlpbytecount0(0)   <= ctlpbytecount(0,0);
ctlpbytecount0(1)   <= ctlpbytecount(0,1);
ctlpbytecount0(2)   <= ctlpbytecount(0,2);
ctlpbytecount0(3)   <= ctlpbytecount(0,3);
ctlpbytecount1(0)   <= ctlpbytecount(1,0);
ctlpbytecount1(1)   <= ctlpbytecount(1,1);
ctlpbytecount1(2)   <= ctlpbytecount(1,2);
ctlpbytecount1(3)   <= ctlpbytecount(1,3);


blk_lnk_up_latch_proc: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         blk_lnk_up_latch <= '1';
         blk_lnk_up_d     <= '0';
      else
         blk_lnk_up_d     <= blk_lnk_up;
         if blk_lnk_up = '0' then
            blk_lnk_up_latch <= '0';
         elsif cpltargetpipeline = ctargetpipeline and blk_lnk_up_latch = '0' then
            blk_lnk_up_latch <= '1';
         end if;
      end if;
   end if;
end process;

blk_lnk_up_latch_o <= blk_lnk_up_latch;

np_req_mode: if C_TRN_NP_FC = "TRUE" generate begin
np_pkt_complete_proc : process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         np_pkt_complete <= (others => '0');
      else
 np_pkt_complete <= rdndreqpipelinedecr & rdreqpipelinedecr;
      end if;
   end if;
end process;

np_pkt_complete_o  <= np_pkt_complete;
end generate;

np_ok_mode: if C_TRN_NP_FC = "FALSE" generate begin
rdndreqpipeline_o  <= rdndreqpipeline;
rdreqpipeline_o    <= rdreqpipeline;
end generate;

data_width_32: if C_S_AXIS_DATA_WIDTH = 32 generate
rd_master_ingress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cr_tready_sig    <= '0';
         rdreqpipelineincr   <= '0';
         rdtargetpipeline    <= (others => '0');
         tlplengthsig        <= (others => '0');
         firstdwbesig        <= (others => '0');
         lastdwbesig         <= (others => '0');
         tlpaddrhigh         <= (others => '0');
         tlpaddrlow          <= (others => '0');
         tlpfmtsig           <= (others => '0');
         rdreqsmsig          <= init;
         rdreq               <= '0';
         badreadreq          <= '0';
         zerolenreadreq      <= '0';
         rdndreqpipelineincr <= '0';
         rdndtargetpipeline  <= "000";
         s_axis_cr_tusersig <= (others => (others => '0'));
         s_axis_cr_tusersigtemp <= (others => '0');
      else
         case rdreqsmsig is
            when init =>
               rdreqpipelineincr <= '0';
               rdndreqpipelineincr <= '0';
               rdreq <= '0';
               if lnkdowndataflush = '0' and blk_lnk_up_latch = '1' then
                  s_axis_cr_tready_sig <= '1';
                  rdreqsmsig       <= memrdreq;
               end if;
            
            when memrdreq =>
               rdreq <= '0';
               rdreqpipelineincr <= '0';
               rdndreqpipelineincr <= '0';
               if blk_lnk_up_latch = '1' then
                  if s_axis_cr_tvalid = '1' then
                     -- Nam - double check
                     -- coverage off -item b 1 -allfalse
                     if s_axis_cr_tdata(30) = '0' then
                        -- Nam - double check
                        -- coverage off -item b 1 -allfalse                     
                        if s_axis_cr_tdata(28 downto 24) = "00000" then
                           -- Nam -- enhance bridge does not foward bad request -- tool issue, work work when the if statement is more than 1 line
                           -- coverage off -item bc 1 -allfalse -condrow 4 5
                           if (s_axis_cr_tuser(2) = '1' or s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or 
                              s_axis_cr_tuser(6) = '1') then
                              badreadreq <= '0';
                           else
                              badreadreq <= '1';
                           end if;
                           tlpattrsig <= s_axis_cr_tdata(13 downto 12);
                           tlpfmtsig    <= s_axis_cr_tdata(30 downto 29);
                           tlplengthsig <= s_axis_cr_tdata(9 downto 0);
                           tlptcsig     <= s_axis_cr_tdata(22 downto 20);
                           rdreqsmsig   <= latch_reqid_tag_be;
                        --else
                        --   rdreqsmsig       <= memrdreq;
                        end if;
                     --else
                     --   rdreqsmsig          <= memrdreq;
                     end if;
                  end if;
                  rdreq <= '0';
               -- Nam - extremely hard to hit case - we covered this in the weekend run with 2 hits
               -- coverage off   
               else
                  --rdtargetpipeline    <= cpltargetpipeline;
                  if s_axis_cr_tvalid = '1' then
                     rdreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            -- Nam - extremely hard to hit, we covered this in the weekend run - 2 hits
            -- coverage off
            when blklinkdown =>
               -- Nam - enhanced bridge doesnot throttle
               -- coverage off -item b 1 -allfalse                       
               if s_axis_cr_tvalid = '1' then
                  if s_axis_cr_tlast = '1' then
                     rdreqsmsig       <= init;
                     s_axis_cr_tready_sig <= '0';
                  end if;
               end if;
            -- coverage on
            when latch_reqid_tag_be =>
               if blk_lnk_up_latch = '1' then
                  -- Nam - enhanced bridge doesnot throttle
                  -- coverage off -item b 1 -allfalse              
                  if s_axis_cr_tvalid = '1' then
                     lastdwbesig  <= s_axis_cr_tdata(7 downto 4);
                     firstdwbesig <= s_axis_cr_tdata(3 downto 0);
                     requesteridsig  <= s_axis_cr_tdata(31 downto 16);
                     tagsig          <= s_axis_cr_tdata(15 downto 8);
                     if tlpfmtsig(0) = '0' then
                        rdreqsmsig  <= latchaddrl;
                     else
                        rdreqsmsig <= latchaddrh;
                     end if;
                     if s_axis_cr_tdata(3 downto 0) = "0000" then
                        zerolenreadreq   <= '1';
                     end if;
                  end if;
               -- Nam - extremely hard to hit case   - we covered this in the weekend run with 2 hits
               -- coverage off                    
               else
                  rdreqsmsig       <= blklinkdown;
               end if;
               -- coverage on
            
            when latchaddrh =>
               if blk_lnk_up_latch = '1' then
                  -- Nam - enhanced bridge doesnot throttle
                  -- coverage off -item b 1 -allfalse   
                  if s_axis_cr_tvalid = '1' then
                     tlpaddrhigh <= s_axis_cr_tdata;
                     rdreqsmsig  <= latchaddrl;
                  end if;
               -- Nam - extremely hard to hit case   
               -- coverage off                    
               else
                  rdreqsmsig       <= blklinkdown;
               end if;
               -- coverage on
            when latchaddrl =>
               if blk_lnk_up_latch = '1' then
                  -- Nam - enhanced bridge doesnot throttle
                  -- coverage off -item bc 1 -allfalse -condrow 1 2               
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     --badreadreq asserted for no bar hit on readreq(root port only)
                     if badreadreq = '0' and zerolenreadreq = '0' then
                        if rdreqpipeline /= "100" then
                           tlpaddrlow <= s_axis_cr_tdata(31 downto 2) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                           tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(31 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(31 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(6 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if conv_integer(tlplengthsig) /= 0 then
                           --when len/=1024DW
                              if conv_integer(tlplengthsig) /= 1 then
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                       firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                             firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                                conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                   lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                       conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                          conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                             firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                                (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                                   firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                                      conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) and 
                                                         firstdwbesig(0)), 12);
                              end if;
                           else
                           --when len=1024DW
                              if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) 
                                       or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                          conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                             firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                                conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                   lastdwbesig(2) or lastdwbesig(3))), 12);
                              -- Nam - extremely hard to hit case   - we covered this in the weekend run with 2 hits
                              -- coverage off                             
                              else
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                              end if;
                              -- coverage on
                           end if;
                           tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= requesteridsig;
                           tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= tagsig;
                           tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= tlptcsig;
                           tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                              blk_function_number;
                           tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpattrsig;
                           tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                           tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                           rdreq <= '1';
                           rdreqsmsig  <= memrdreq;
                           rdreqpipelineincr <= '1';
                           rdtargetpipeline <= rdtargetpipeline + 1;
                           if (orrdreqpipeline /= rdtargetpipeline) and
                           (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                              wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                           else
                              wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                           end if;
                           if C_PCIEBAR_AS = 0 then
                              s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(C_PCIEBAR_NUM-1 downto 0) <= 
                                 s_axis_cr_tuser(C_PCIEBAR_NUM+1 downto 2);
                           else
                              for i in 0 to C_PCIEBAR_NUM-1 loop
                                 s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(i) <= s_axis_cr_tuser(2*(i+1));
                              end loop;
                           end if;
                        else
                           s_axis_cr_tready_sig <= '0';
                           rdreqsmsig   <= throttle;
                           tlpaddrlow <= s_axis_cr_tdata(31 downto 2) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if C_PCIEBAR_AS = 0 then
                              s_axis_cr_tusersigtemp(C_PCIEBAR_NUM-1 downto 0) <= s_axis_cr_tuser(C_PCIEBAR_NUM+1 downto 2);
                           else
                              for i in 0 to C_PCIEBAR_NUM-1 loop
                                 s_axis_cr_tusersigtemp(i) <= s_axis_cr_tuser(2*(i+1));
                              end loop;
                           end if;
                        end if;
                     else --zero length read for EP/RC also nobarhit for RC
                        if rdndreqpipeline /= "100" then
                           rdreqsmsig  <= memrdreq;
                           if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend or 
                             badreadreq = '1' then
                              wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                           else
                              wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                           end if;
                           tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlptcsig;
                           tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlpattrsig;
                           tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= requesteridsig;
                           tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                              blk_function_number;
                           tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= tagsig;
                           rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(6 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                 conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if badreadreq = '1' then
                              cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                           elsif zerolenreadreq = '1' then
                              cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                           end if;
                           rdndtargetpipeline <= rdndtargetpipeline +1;
                           rdndreqpipelineincr <= '1';
                           badreadreq <= '0';
                           zerolenreadreq <= '0';
                           -- NAM / JRH Tool bug doesn't exclude the second condition. removed cov off item b 2. Moved cov off.
                           if conv_integer(tlplengthsig) /= 0 then
                           --when len/=1024DW
                              -- coverage off -item b 1
                              if conv_integer(tlplengthsig) /= 1 then
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                       firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                       conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                          conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                             firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                                (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                                   firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                                      conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) 
                                                         and firstdwbesig(0)), 12);
                              end if;
                           -- NAM / JRH Tool bug doesn't exclude the second condition. Moved cov off.
                           else
                           --when len=1024DW
                              if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) 
                                       or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                          conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                             firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) 
                                                + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                   lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                              end if;
                           end if;
                        else
                           s_axis_cr_tready_sig <= '0';
                           rdreqsmsig   <= throttle_nd;
                           rdndtlpaddrlow <= 
                              s_axis_cr_tdata(6 downto 2) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                        end if; 
                     end if;
                  end if;
               -- Nam - extremely hard to hit case - we covered this in the weekend run with 2 hits
               -- coverage off                    
               else
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     rdreqsmsig       <= init;
                     s_axis_cr_tready_sig <= '0';
                  else
                     rdreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            
            when throttle =>
               if blk_lnk_up_latch = '1' then
                  if rdreqpipeline /= "100" then
                    --pipeline full for CplD (i.e., compl with data)
                     tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0)))    <= tlpaddrlow;
                     tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0)))    <= tlpaddrlow;
                     rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpaddrlow(6 downto 0);
                     if conv_integer(tlplengthsig) /= 0 then
                     --when len/=1024DW
                        if conv_integer(tlplengthsig) /= 1 then
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                 firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                    conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                       conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                          firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                             conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                 conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + conv_integer(not((firstdwbesig(3) 
                                    xor firstdwbesig(1)) or (firstdwbesig(2) xor firstdwbesig(0)))) + conv_integer((firstdwbesig(3)
                                       and firstdwbesig(0)) and (firstdwbesig(2) nor firstdwbesig(1))) + 
                                          conv_integer((firstdwbesig(3) and firstdwbesig(0)) and (firstdwbesig(2) nand 
                                             firstdwbesig(1))) - conv_integer(firstdwbesig(3) and firstdwbesig(2) and 
                                                firstdwbesig(1) and firstdwbesig(0)), 12);
                        end if;
                     else
                     --when len=1024DW
                        if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + conv_integer(firstdwbesig(2) 
                                    or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(2) or lastdwbesig(3)) + 
                                       conv_integer(firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(1) or 
                                          lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(0) or lastdwbesig(1) or lastdwbesig(2) or 
                                                lastdwbesig(3))), 12);
                        -- Nam - extremely hard to hit case - we covered this in the weekend run with 6 hits
                        -- coverage off                                                    
                        else
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                        end if;
                        -- coverage on
                     end if;
                     tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= requesteridsig;
                     tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= tagsig;
                     tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= tlptcsig;
                     tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                        blk_function_number;
                     tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpattrsig;
                     tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                     tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                     rdreq <= '1';
                     --if blk_lnk_up = '0' then
                     --   s_axis_cr_tready_sig <= '0';
                     --   rdreqsmsig  <= init;
                     --else
                     rdreqsmsig  <= memrdreq;
                     s_axis_cr_tready_sig <= '1';
                     --end if;
                     rdreqpipelineincr <= '1';
                     rdtargetpipeline <= rdtargetpipeline + 1;
                     if (orrdreqpipeline /= rdtargetpipeline) and
                     (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                        wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                     else
                        wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                     end if;
                     s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tusersigtemp;
                  end if;
               else
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
               end if;
            
            when throttle_nd =>
               if blk_lnk_up_latch = '1' then
                  if rdndreqpipeline /= "100" then
                    --pipeline full for Cpl (i.e., compl without data - no barhit or zero len)
                     --if blk_lnk_up = '0' then
                     --   s_axis_cr_tready_sig <= '0';
                     --   rdreqsmsig  <= init;
                     --else
                     rdreqsmsig  <= memrdreq;
                     s_axis_cr_tready_sig <= '1';
                     --end if;
                     if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend or 
                       badreadreq = '1' then
                        wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                     else
                        wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                     end if;
                     tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlptcsig;
                     tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlpattrsig;
                     tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= requesteridsig;
                     tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                        blk_function_number;
                     tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= tagsig;
                     rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= rdndtlpaddrlow;
                     if badreadreq = '1' then
                        cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                     elsif zerolenreadreq = '1' then
                        cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                     end if;
                     rdndtargetpipeline <= rdndtargetpipeline +1;
                     rdndreqpipelineincr <= '1';
                     badreadreq <= '0';
                     zerolenreadreq <= '0';
                     -- NAM / JRH Tool bug doesn't exclude the second condition. removed cov off item b 2. Moved cov off.
                     if conv_integer(tlplengthsig) /= 0 then
                     --when len/=1024DW
                        -- coverage off -item b 1
                        if conv_integer(tlplengthsig) /= 1 then
                           -- Not hit for EP, include for RC
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                 firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                    conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                       conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                          firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                             conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                 conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + conv_integer(not((firstdwbesig(3) 
                                    xor firstdwbesig(1)) or (firstdwbesig(2) xor firstdwbesig(0)))) + conv_integer((firstdwbesig(3)
                                       and firstdwbesig(0)) and (firstdwbesig(2) nor firstdwbesig(1))) + 
                                          conv_integer((firstdwbesig(3) and firstdwbesig(0)) and (firstdwbesig(2) nand 
                                             firstdwbesig(1))) - conv_integer(firstdwbesig(3) and firstdwbesig(2) and 
                                                firstdwbesig(1) and firstdwbesig(0)), 12);
                        end if;
                     -- NAM / JRH Tool bug doesn't exclude the second condition. Moved cov off.
                     -- coverage off
                     else
                     --when len=1024DW
                           -- Not hit for EP, include for RC
                        if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + conv_integer(firstdwbesig(2) 
                                    or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(2) or lastdwbesig(3)) + 
                                       conv_integer(firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(1) or 
                                          lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(0) or lastdwbesig(1) or lastdwbesig(2) or 
                                                lastdwbesig(3))), 12);
                        else
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                        end if;
                           -- coverage on
                     end if;
                  end if;
               -- Nam - extremely hard to hit cases - requires zero length request right at link_down
               -- coverage off                    
               else
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
               end if;
               -- coverage on
            
            -- coverage off
            when others => 
               rdreqsmsig <= init;
            -- coverage on
         end case;
         if blk_lnk_up_latch = '0' and cpltargetpipeline /= ctargetpipeline then
            rdtargetpipeline <= addrstreampipeline;
         end if;
      end if;
   end if;
end process;

cplnd_master_egress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         cplndtlpsmsig <= memcplcrtdatabeat1;
         cplndtargetpipeline <= "000";
         rdndreqpipelinedecr <= '0';
         m_axis_cc_tvalid_nd <= '0';
         m_axis_cc_tdata_nd <= (others => '0');
         m_axis_cc_tstrb_nd <= (others => '0');
         m_axis_cc_tlast_nd <= '0';
         dis_valid_nd <= '0';
         orcplndpipeline <= (others => '0');
         cplndpendcpl <= (others => '0');
      else
         if orcplndpipeline /= rdndtargetpipeline then
            cplndpendcpl(conv_integer(orcplndpipeline(1 downto 0))) <= '0';
            if master_wr_idle = '1' or wrpendflush(conv_integer(orcplndpipeline(1 downto 0)))(2 downto 0) = wrreqcomp
                       or wrpendflush(conv_integer(orcplndpipeline(1 downto 0)))(3) = '1' then
               cplndpendcpl(conv_integer(orcplndpipeline(1 downto 0))) <= '1';
               orcplndpipeline <= orcplndpipeline + 1;
            end if;
         end if;
        
         -- cplndpendcpl needs to be reset on link down event
         if blk_lnk_up_latch = '0' then
            cplndpendcpl <= (others => '0');
         end if;
         case cplndtlpsmsig is
            when memcplcrtdatabeat1 =>
               rdndreqpipelinedecr <= '0';
               m_axis_cc_tvalid_nd <= '0';
               m_axis_cc_tlast_nd <= '0';
               m_axis_cc_tstrb_nd <= x"0";
               if cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline then
                  if blk_lnk_up_latch = '1' then
                     if cplndpendcpl(conv_integer(cplndtargetpipeline(1 downto 0))) = '1' then
                        if cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) = "000" then
                          m_axis_cc_tdata_nd <= '0' & "10" & "01010" & '0' & tlpndtc(conv_integer(cplndtargetpipeline(1 downto 0)))
                            & "0000" & '0' & '0' & tlpndattr(conv_integer(cplndtargetpipeline(1 downto 0))) & "00" & "0000000001";
                        -- coverage off
                        else
                          m_axis_cc_tdata_nd <= '0' & "00" & "01010" & '0' & tlpndtc(conv_integer(cplndtargetpipeline(1 downto 0)))
                             & "0000" & '0' & '0' & tlpndattr(conv_integer(cplndtargetpipeline(1 downto 0))) & "00" & "0000000000";
                        -- coverage on
                        end if;
                        m_axis_cc_tstrb_nd <= (others => '1');
                        m_axis_cc_tvalid_nd <= '1';
                        if m_axis_cc_tready = '1' and m_axis_cc_tvalid_nd = '1' then
                           cplndtlpsmsig <= memcplcrtdatabeat2;
                           if cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) = "000" then
                              m_axis_cc_tdata_nd <= tlpndcompleterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                 cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & x"001";
                           -- coverage off
                           else
                              m_axis_cc_tdata_nd <= tlpndcompleterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                 cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                                    tlpndbytecount(conv_integer(cplndtargetpipeline(1 downto 0)));
                           -- coverage on
                           end if;
                        --else
                        --   cplndtlpsmsig <= memcplcrtdatabeat1;
                        end if;
                     end if;
                  -- Nam - extremely hard to hit cases   
                  -- coverage off                       
                  else
                     cplndtlpsmsig       <= memcplcrtdatabeat1;
                     rdndreqpipelinedecr <= '1';
                     cplndtargetpipeline <= cplndtargetpipeline + 1;
                  end if;
                  -- coverage on
               end if;
            
            when memcplcrtdatabeat2 =>
               m_axis_cc_tstrb_nd <= (others => '1');
               m_axis_cc_tvalid_nd <= '1';
               -- Nam - enhanced bridge doesnot throttle
               -- coverage off -item bc 1 -allfalse -condrow 2 3               
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tdata_nd <= tlpndrequesterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                     tlpndtag(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                        rdndtlpaddrl(conv_integer(cplndtargetpipeline(1 downto 0)));
                  if cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) = "000" then
                     cplndtlpsmsig <= memcplcrtdatabeat3;
                  -- coverage off
                  else
                     cplndtlpsmsig <= transfer_complete;
                     m_axis_cc_tlast_nd <= '1';
                  -- coverage on
                  end if;
               --else
               --   cplndtlpsmsig <= memcplcrtdatabeat2;
               end if;
            
            when memcplcrtdatabeat3 =>
               m_axis_cc_tstrb_nd <= (others => '1');
               m_axis_cc_tvalid_nd <= '1';
               -- Nam - enhanced bridge doesnot throttle
               -- coverage off -item b 1 -allfalse
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tdata_nd <= x"00000000";
                  m_axis_cc_tlast_nd <= '1';
                  cplndtlpsmsig <= transfer_complete;
               --else
               --   cplndtlpsmsig <= memcplcrtdatabeat3;
               end if;
            
            when transfer_complete =>
                  if m_axis_cc_tready = '1' then
                  cplndtlpsmsig <= memcplcrtdatabeat1;
                  m_axis_cc_tvalid_nd <= '0';
                  m_axis_cc_tlast_nd <= '0';
                  m_axis_cc_tstrb_nd <= x"0";
                  rdndreqpipelinedecr <= '1';
                  cplndtargetpipeline <= cplndtargetpipeline + 1;
                  end if;

         -- coverage off
         when others =>
            cplndtlpsmsig <= memcplcrtdatabeat1;
         -- coverage on
      end case;
      end if;
   end if;
end process;

cpl_master_egress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         cpltlpsmsig <= memcplpipeline;
         cpltargetpipeline <= (others => '0');
         rdreqpipelinedecr <= '0';
         cplpacket1 <= '0';
         firstdwen   <= '0';
         lnkdowndataflush <= '0';
         m_axis_cc_tvalid_d <= '0';
         m_axis_cc_tstrb_d <= (others => '0');
         m_axis_cc_tlast_d <= '0';
         rd_en_sig <= '0';
         cplcounter <= (others => '0');
         cpldsplitcounttemp <= (others => '0');
         rdtlpaddrltemp <= (others => '0');
         ctlpbytecounttemp <= (others => '0');
         ctlplengthtemp <= (others => '0');
         tlplengthcntr <= (others => '0');
         dis_valid_d <= '0';
         m_axis_cc_tdata_h <= (others => '0');
         data_phase <= '0';
         dis_rden <= '0';
         corruptdataflush <= '0';
         wait_till_not_empty <= '0';
         totallength <= (others => '0');
         totalbytecount <= (others => '0');
         linkdownflushdepth <= (others => '0');
         rrespdelayed <= '0';
      else
         case cpltlpsmsig is
            when memcplpipeline =>
               rdreqpipelinedecr <= '0';
               m_axis_cc_tlast_d <= '0';
               m_axis_cc_tvalid_d <= '0';
               m_axis_cc_tstrb_d <= x"0";
               if blk_lnk_up_latch = '1' then
                  if cplndtargetpipeline = rdndtargetpipeline then
                     if cpltargetpipeline /= ctargetpipeline then
                     --pending completions exist
                        cplcounter <= "00000";
                        cpldsplitcounttemp <= cpldsplitcount(conv_integer(cpltargetpipeline(1 downto 0)));
                        rdtlpaddrltemp <= rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)));
                        ctlpbytecounttemp <= ctlpbytecount0(conv_integer(cpltargetpipeline(1 downto 0)));
                        ctlplengthtemp <= ctlplength0(conv_integer(cpltargetpipeline(1 downto 0)));
                        totallength <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                        linkdownflushdepth <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                        totalbytecount <= tlpbytecount(conv_integer(cpltargetpipeline(1 downto 0)));
                        cplpacket1 <= '1';
                        cpltlpsmsig <= memcplcrtdatabeat1;
                        rrespdelayed <= '0';
                     else
                        cpltlpsmsig <= memcplpipeline;
                     end if;
                  end if;
               elsif cpltargetpipeline /= ctargetpipeline and empty = '0' then
                  cpltlpsmsig <= blklinkdown_corruptdata;
                  lnkdowndataflush <= '1';
                  tlplengthcntr <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                  rd_en_sig <= '1';
               end if;
            
            
            when memcplcrtdatabeat1 =>
               m_axis_cc_tlast_d <= '0';
               rrespdelayed <= rresp(conv_integer(cpltargetpipeline(1 downto 0)))(2);
                  if (((cplpendcpl(conv_integer(cpltargetpipeline(1 downto 0))) = '1' and rrespdelayed = '1') or 
                     slv_write_idle = '1') and rresp(conv_integer(cpltargetpipeline(1 downto 0)))(2) = '1')
                     or blk_lnk_up_latch = '0' then
                  --ordering & rresp check
                     if rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1 downto 0) = "00" then
                     --OKAY response
                        if blk_lnk_up_latch = '1' then
                        --link up
                           m_axis_cc_tdata_h <= '0' & "10" & "01010" & '0' & tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              "0000" & '0' & '0' & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & 
                                              ctlplengthtemp;
                           tlplengthcntr <= ctlplengthtemp;
                           m_axis_cc_tstrb_d <= (others => '1');
                           m_axis_cc_tvalid_d <= '1';
                           if m_axis_cc_tready = '1' and m_axis_cc_tvalid_d = '1' then
                              linkdownflushdepth <= linkdownflushdepth - ctlplengthtemp;
                              cpltlpsmsig <= memcplcrtdatabeat2;
                              m_axis_cc_tdata_h <= tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                 rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & 
                                    '0' & (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                    rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & ctlpbytecounttemp;
                           --else
                           --   cpltlpsmsig <= memcplcrtdatabeat1;
                           end if;
                        else
                        --link is down
                           if empty = '0' then
                              cpltlpsmsig       <= blklinkdown_corruptdata;
                              m_axis_cc_tvalid_d <= '0';
                              tlplengthcntr <= linkdownflushdepth;
                              rd_en_sig            <= '1';
                              lnkdowndataflush <= '1';
                           else
                              cpltlpsmsig       <= memcplpipeline;
                           end if;
                        end if;
                     else
                     --DECERR or SLVERR response
                        if blk_lnk_up_latch = '1' then
                           m_axis_cc_tdata_h <= '0' & "00" & "01010" & '0' & tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              "0000" & '0' & '0' & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & totallength;
                           tlplengthcntr <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                           m_axis_cc_tstrb_d <= (others => '1');
                           m_axis_cc_tvalid_d <= '1';
                           -- Nam - enhanced bridge doesnot throttle
                           -- coverage off -item c 1 -condrow 2
                           if m_axis_cc_tready = '1' and m_axis_cc_tvalid_d = '1' then
                              cpltlpsmsig <= memcplcrtdatabeat2;
                              m_axis_cc_tdata_h <= tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                 rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) &
                                 '0' & (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                    rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & totalbytecount;
                           --else
                           --   cpltlpsmsig <= memcplcrtdatabeat1;
                           end if;
                        -- Nam - extremely hard to hit cases - DECERR or SLVERR with link_down
                        -- coverage off                             
                        else
                           if empty = '0' then
                              cpltlpsmsig       <= blklinkdown_corruptdata;
                              m_axis_cc_tvalid_d <= '0';
                              tlplengthcntr <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                              rd_en_sig            <= '1';
                              lnkdowndataflush <= '1';
                           else
                              cpltlpsmsig       <= memcplpipeline;
                           end if;
                        end if;
                        -- coverage on
                     end if;
                  end if;
            
            when blklinkdown_corruptdata =>
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tvalid_d <= '0';
               end if;
               rdreqpipelinedecr <= '0';
               if empty = '0' then
                  wait_till_not_empty <= '1';
                  if tlplengthcntr /= "0000000001" then
                     tlplengthcntr <= tlplengthcntr - 1;
                     rd_en_sig <= '1';
                  else
                     if lnkdowndataflush = '1' then
                        if cpltargetpipeline + 1 /= ctargetpipeline then
                           tlplengthcntr <= tlplength(conv_integer(cpltargetpipeline(1 downto 0) + 1));
                           --rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                        else
                           -- Nam - enhanced bridge doesnot throttle
                           -- coverage off -item bc 1 -allfalse -condrow 2 3
                           if m_axis_cc_tvalid_d = '0' or m_axis_cc_tready = '1' then
                              cpltlpsmsig <= memcplpipeline;
                              --rdreqpipelinedecr <= '1';
                              cpltargetpipeline <= cpltargetpipeline + 1;
                              wait_till_not_empty <= '0';
                           end if;
                           rd_en_sig <= '0';
                           lnkdowndataflush <= '0';
                        end if;
                     else
                        -- Nam - enhanced bridge doesnot throttle
                        -- coverage off -item bc 1 -allfalse -condrow 2 3                  
                        if m_axis_cc_tvalid_d = '0' or m_axis_cc_tready = '1' then
                           cpltlpsmsig <= memcplpipeline;
                           rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                           wait_till_not_empty <= '0';
                        end if;
                        rd_en_sig <= '0';
                        corruptdataflush <= '0';
                     end if;
                  end if;
               end if;

            when memcplcrtdatabeat2 =>
               if rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1 downto 0) = "00" then
                  m_axis_cc_tstrb_d <= (others => '1');
                  m_axis_cc_tvalid_d <= '1';
                  -- Nam - enhanced bridge doesnot throttle
                  -- coverage off -item b 1 -allfalse
                  if m_axis_cc_tready = '1' then
                     if cplpacket1 <= '0' then
                        m_axis_cc_tdata_h <= tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                           tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & x"00";
                     else
                        m_axis_cc_tdata_h <= tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                           tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp;
                     end if;
                     cpltlpsmsig <= memcpltxdata;
                     firstdwen   <= '1';
                  --else
                  --   cpltlpsmsig <= memcplcrtdatabeat2;
                  end if;
               else
                  m_axis_cc_tstrb_d <= (others => '1');
                  m_axis_cc_tvalid_d <= '1';
                  -- Nam - enhanced bridge doesnot throttle
                  -- coverage off -item b 1 -allfalse
                  if m_axis_cc_tready = '1' then
                     m_axis_cc_tdata_h <= tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                        tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp;
                     m_axis_cc_tlast_d <= '1';
                     cpltlpsmsig <= blklinkdown_corruptdata;
                     tlplengthcntr <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                     rd_en_sig <= '1';
                     corruptdataflush <= '1';
                  --else
                  --   cpltlpsmsig <= memcplcrtdatabeat2;
                  end if;
               end if;
            
            when memcpltxdata =>
               if empty = '0' or tlplengthcntr = "0000000000" then
                  -- Nam - enhanced bridge doesnot throttle
                  -- coverage off -item b 1 -allfalse
                  if m_axis_cc_tready = '1' then
                     m_axis_cc_tvalid_d <= not(empty);
                     data_phase <= '1';
                     if tlplengthcntr = "0000000001" then
                        m_axis_cc_tlast_d <= '1';
                     end if;
                     if firstdwen = '1' then
                        m_axis_cc_tstrb_d <= x"F";
                        firstdwen <= '0';
                        tlplengthcntr <= tlplengthcntr - 1;
                     elsif tlplengthcntr = "0000000000" then
                        m_axis_cc_tlast_d <= '0';
                        data_phase <= '0';
                        m_axis_cc_tvalid_d <= '0';
                        if cplcounter /= cpldsplitcounttemp then
                           cpltlpsmsig <= memcplcrtdatabeat1;
                           cplcounter <= cplcounter + 1;
                           if cplcounter /= "00000" then
                              ctlpbytecounttemp <= ctlpbytecounttemp - 
                                 (ctlplength1(conv_integer(cpltargetpipeline(1 downto 0))) & "00");
                           else
                              ctlpbytecounttemp <= ctlpbytecounttemp - 
                                 ctlpbytecount1(conv_integer(cpltargetpipeline(1 downto 0)));
                           end if;
                           if cplcounter+1 /= cpldsplitcounttemp then
                              ctlplengthtemp <= ctlplength1(conv_integer(cpltargetpipeline(1 downto 0)));
                           else
                              ctlplengthtemp <= ctlplength2(conv_integer(cpltargetpipeline(1 downto 0)));
                           end if;
                           cplpacket1 <= '0';
                        else
                           m_axis_cc_tstrb_d <= x"F";
                           cpltlpsmsig <= memcplpipeline;
                           rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                        end if;
                     else
                        m_axis_cc_tstrb_d <= (others => '1');
                        tlplengthcntr <= tlplengthcntr - 1;
                     end if;
                  end if;
               end if;
         
         -- coverage off
            when others =>
            cpltlpsmsig <= memcplpipeline;
         -- coverage on
         end case;
         --if blk_lnk_up = '0' and blk_lnk_up_d = '1' then
            --cpltargetpipeline <= cpltargetpipeline - rdreqpipeline;
         --end if;
      end if;
   end if;
end process;
end generate;

data_width_64: if C_S_AXIS_DATA_WIDTH = 64 generate
rd_master_ingress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cr_tready_sig    <= '0';
         rdreqpipelineincr   <= '0';
         rdtargetpipeline    <= (others => '0');
         tlplengthsig        <= (others => '0');
         firstdwbesig        <= (others => '0');
         lastdwbesig         <= (others => '0');
         tlpaddrhigh         <= (others => '0');
         tlpaddrlow          <= (others => '0');
         tlpfmtsig           <= (others => '0');
         rdreqsmsig          <= init;
         rdreq               <= '0';
         badreadreq          <= '0';
         zerolenreadreq      <= '0';
         rdndreqpipelineincr <= '0';
         rdndtargetpipeline  <= "000";
         s_axis_cr_tusersig <= (others => (others => '0'));
         s_axis_cr_tusersigtemp <= (others => '0');
      else
         case rdreqsmsig is
            when init =>
               rdreqpipelineincr <= '0';
               rdndreqpipelineincr <= '0';
               rdreq <= '0';
               if lnkdowndataflush = '0' and blk_lnk_up_latch = '1' then
                  s_axis_cr_tready_sig <= '1';
                  rdreqsmsig       <= memrdreq;
               end if;
            
            when memrdreq =>
               rdreq <= '0';
               if blk_lnk_up_latch = '1' then
                  if s_axis_cr_tvalid = '1' then
                     -- Nam - double check, bit 30 always = 0
                     -- coverage off -item b 1 -allfalse                  
                     if s_axis_cr_tdata(30) = '0' then
                        -- Nam - core does not support mem read locked
                        -- coverage off -item b 1 -allfalse
                        if s_axis_cr_tdata(28 downto 24) = "00000" then
                           -- Nam - enhance bridge does not forward bad request -- tool issue, work work when the if statement is more than 1 line
                           -- coverage off -item bc 1 -allfalse -condrow 5
                           if ((s_axis_cr_tuser(2) = '1' and C_PCIEBAR_NUM = 1) or (C_PCIEBAR_NUM > 1 and (s_axis_cr_tuser(2) = '1' or 
                             s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) then
                              badreadreq <= '0';
                           else
                              badreadreq <= '1';
                           end if;
                              tlpattrsig <= s_axis_cr_tdata(13 downto 12);
                              tlpfmtsig    <= s_axis_cr_tdata(30 downto 29);
                              tlplengthsig <= s_axis_cr_tdata(9 downto 0);
                              tlptcsig     <= s_axis_cr_tdata(22 downto 20);
                              lastdwbesig  <= s_axis_cr_tdata(39 downto 36);
                              firstdwbesig <= s_axis_cr_tdata(35 downto 32);
                              requesteridsig  <= s_axis_cr_tdata(63 downto 48);
                              tagsig          <= s_axis_cr_tdata(47 downto 40);
                                 if s_axis_cr_tdata(29) = '0' then
                                    rdreqsmsig  <= latchaddrl;
                                 else
                                    rdreqsmsig <= latchaddrh;
                                 end if;
                              if s_axis_cr_tdata(35 downto 32) = "0000" then
                                 zerolenreadreq   <= '1';
                              end if;
                        --else
                        --   rdreqsmsig       <= memrdreq;
                        end if;
                     --else
                     --   rdreqsmsig          <= memrdreq;
                     end if;
                  end if;
                  rdreq <= '0';
               -- Nam - extremely hard to hit case
               -- coverage off                      
               else
                  --rdtargetpipeline    <= cpltargetpipeline;
                  if s_axis_cr_tvalid = '1' then
                     rdreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
               rdreqpipelineincr <= '0';
               rdndreqpipelineincr <= '0';
            
            -- Nam - extremely hard to hit case
            -- coverage off    
            when blklinkdown =>
               if s_axis_cr_tvalid = '1' then
                  if s_axis_cr_tlast = '1' then
                     rdreqsmsig       <= init;
                     s_axis_cr_tready_sig <= '0';
                  end if;
               end if;
            -- coverage on
            
            when latchaddrh =>
               if blk_lnk_up_latch = '1' then
                  -- Nam - enhanced bridge doesn't throttle
                  -- coverage off -item bc 1 -condrow 1
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     -- Nam - never hit condition
                     -- coverage off -item c 1 -condrow 1 2
                     if badreadreq = '0' and zerolenreadreq = '0' then
                        if rdreqpipeline /= "100" then
                           tlpaddrlow <= s_axis_cr_tdata(63 downto 34) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) +
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                           tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(63 downto 34) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(63 downto 34) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(38 downto 34) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if conv_integer(tlplengthsig) /= 0 then
                           --when len/=1024DW
                              if conv_integer(tlplengthsig) /= 1 then
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                       firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                       conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                          conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                             firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                                (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                                   firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                                      conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) and 
                                                         firstdwbesig(0)), 12);
                              end if;
                           else
                           --when len=1024DW
                              if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) 
                                       or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                                                      
                              -- Nam - extremely hard to hit case - we covered this in the weekend run with 1 hits
                              -- coverage off                                  
                              else
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                              end if;
                              -- coverage on
                           end if;
                           tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= requesteridsig;
                           tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= tagsig;
                           tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= tlptcsig;
                           tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                              blk_function_number;
                           tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpattrsig;
                           tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                           tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                           rdreq <= '1';
                           rdreqsmsig  <= memrdreq;
                           rdreqpipelineincr <= '1';
                           rdtargetpipeline <= rdtargetpipeline + 1;
                           if (orrdreqpipeline /= rdtargetpipeline) and
                           (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                              wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                           else
                              wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                           end if;
                           for i in 0 to C_PCIEBAR_NUM-1 loop
                              s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(i) <= s_axis_cr_tuser(2*(i+1));
                           end loop;
                        else
                           s_axis_cr_tready_sig <= '0';
                           rdreqsmsig   <= throttle;
                           tlpaddrlow <= s_axis_cr_tdata(63 downto 34) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) +
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                           for i in 0 to C_PCIEBAR_NUM-1 loop
                              s_axis_cr_tusersigtemp(i) <= s_axis_cr_tuser(2*(i+1));
                           end loop;
                        end if;
                     else
                        if rdndreqpipeline /= "100" then
                           rdreqsmsig  <= memrdreq;
                           if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend or 
                             badreadreq = '1' then
                              wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                           else
                              wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                           end if;
                           tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlptcsig;
                           tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlpattrsig;
                           tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= requesteridsig;
                           tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                              blk_function_number;
                           tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= tagsig;
                           rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(38 downto 34) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if badreadreq = '1' then
                              cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                           elsif zerolenreadreq = '1' then
                              cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                           end if;
                           rdndtargetpipeline <= rdndtargetpipeline +1;
                           rdndreqpipelineincr <= '1';
                           badreadreq <= '0';
                           zerolenreadreq <= '0';
                           -- NAM / JRH Tool bug doesn't exclude the second condition. removed cov off item b 2. Moved cov off.
                           if conv_integer(tlplengthsig) /= 0 then
                           --when len/=1024DW
                              -- coverage off -item b 1
                              if conv_integer(tlplengthsig) /= 1 then
                           -- Not hit for EP, include for RC
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                       firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                       conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                          conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                             firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                                (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                                   firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                                      conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) and 
                                                         firstdwbesig(0)), 12);
                              end if;
                           -- NAM / JRH Tool bug doesn't exclude the second condition. Moved cov off.
                           -- coverage off
                           else
                           --when len=1024DW
                           -- Not hit for EP, include for RC
                              if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) 
                                       or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                       conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                          conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                             firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                                conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                   lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                              end if;
                           -- coverage on
                           end if;
                        else
                           s_axis_cr_tready_sig <= '0';
                           rdreqsmsig   <= throttle_nd;
                           rdndtlpaddrlow <= 
                              s_axis_cr_tdata(38 downto 34) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                        end if;
                     end if;
                  end if;
               
               -- Nam - extremely hard to hit case - we covered this in the weekend run with 2 hits
               -- coverage off                      
               else
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     rdreqsmsig       <= init;
                     s_axis_cr_tready_sig <= '0';
                  else
                     rdreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
               
            when latchaddrl =>
               if blk_lnk_up_latch = '1' then
                  -- Nam - enhance bridge doesn't throttle
                  -- coverage off -item bc 1 -allfalse -condrow 1 2
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     -- Nam - never hit condition
                     -- coverage off -item c 1 -condrow 1
                     if badreadreq = '0' and zerolenreadreq = '0' then
                        if rdreqpipeline /= "100" then
                           tlpaddrlow <= s_axis_cr_tdata(31 downto 2) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                           tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(31 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(31 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(6 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if conv_integer(tlplengthsig) /= 0 then
                           --when len/=1024DW
                              if conv_integer(tlplengthsig) /= 1 then
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                       firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))
                                                  + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                     or lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                       conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                          conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                             firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                                (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                                   firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                                      conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) and 
                                                         firstdwbesig(0)), 12);
                              end if;
                           else
                           --when len=1024DW
                              if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) 
                                       or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                                                      
                              -- Nam - extremely hard to hit case - we covered this in the weekend run with 4 hits
                              -- coverage off                                                          
                              else
                                 tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                              end if;
                              -- coverage on
                           end if;
                           tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= requesteridsig;
                           tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= tagsig;
                           tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= tlptcsig;
                           tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                              blk_function_number;
                           tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpattrsig;
                           tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                           tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                           rdreq <= '1';
                           rdreqsmsig  <= memrdreq;
                           rdreqpipelineincr <= '1';
                           rdtargetpipeline <= rdtargetpipeline + 1;
                           if (orrdreqpipeline /= rdtargetpipeline) and
                           (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                              wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                           else
                              wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                           end if;
                           if C_PCIEBAR_AS = 0 then
                              s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(C_PCIEBAR_NUM-1 downto 0) <= 
                                 s_axis_cr_tuser(C_PCIEBAR_NUM+1 downto 2);
                           else
                              for i in 0 to C_PCIEBAR_NUM-1 loop
                                 s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(i) <= s_axis_cr_tuser(2*(i+1));
                              end loop;
                           end if;
                        else
                           s_axis_cr_tready_sig <= '0';
                           rdreqsmsig   <= throttle;
                           tlpaddrlow <= s_axis_cr_tdata(31 downto 2) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                              conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if C_PCIEBAR_AS = 0 then
                              s_axis_cr_tusersigtemp(C_PCIEBAR_NUM-1 downto 0) <= s_axis_cr_tuser(C_PCIEBAR_NUM+1 downto 2);
                           else
                              for i in 0 to C_PCIEBAR_NUM-1 loop
                                 s_axis_cr_tusersigtemp(i) <= s_axis_cr_tuser(2*(i+1));
                              end loop;
                           end if;
                        end if;
                     else
                        if rdndreqpipeline /= "100" then
                           rdreqsmsig  <= memrdreq;
                           if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend or 
                             badreadreq = '1' then
                              wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                           else
                              wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                           end if;
                           tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlptcsig;
                           tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlpattrsig;
                           tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= requesteridsig;
                           tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                              blk_function_number;
                           tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= tagsig;
                           rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(6 downto 2) & 
                              conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + conv_integer(not(firstdwbesig(1) or 
                                 firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0))) + 
                                   conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)))), 2);
                           if badreadreq = '1' then
                              cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                           elsif zerolenreadreq = '1' then
                              cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                           end if;
                           rdndtargetpipeline <= rdndtargetpipeline +1;
                           rdndreqpipelineincr <= '1';
                           badreadreq <= '0';
                           zerolenreadreq <= '0';
                           -- coverage off
                           if conv_integer(tlplengthsig) /= 0 then
                           --when len/=1024DW
                              if conv_integer(tlplengthsig) /= 1 then
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                       firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) 
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                           -- coverage on
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                       conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                          conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                             firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                                (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                                   firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                                      conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) and 
                                                         firstdwbesig(0)), 12);
                           -- coverage off
                              end if;
                           else
                           --when len=1024DW
                              if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                    conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or
                                       firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                          conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                                firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) 
                                                   + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) 
                                                      or lastdwbesig(2) or lastdwbesig(3))), 12);
                              else
                                 tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                              end if;
                           end if;
                           -- coverage on
                        else
                           s_axis_cr_tready_sig <= '0';
                           rdreqsmsig   <= throttle_nd;
                           rdndtlpaddrlow <= 
                              s_axis_cr_tdata(6 downto 2) & conv_std_logic_vector((conv_integer(not(firstdwbesig(0))) + 
                                 conv_integer(not(firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(2) or 
                                    firstdwbesig(1) or firstdwbesig(0))) + conv_integer(not(firstdwbesig(3) or firstdwbesig(2) or 
                                       firstdwbesig(1) or firstdwbesig(0)))), 2);
                        end if;
                     end if;
                  end if;

               -- Nam - extremely hard to hit case
               -- coverage off                      
               else
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     rdreqsmsig       <= init;
                     s_axis_cr_tready_sig <= '0';
                  else
                     rdreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            
            when throttle =>
               if blk_lnk_up_latch = '1' then
                  if rdreqpipeline /= "100" then
                    --pipeline full for CplD (i.e., compl with data)
                     tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0)))    <= tlpaddrlow;
                     tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0)))    <= tlpaddrlow;
                     rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpaddrlow(6 downto 0);
                     if conv_integer(tlplengthsig) /= 0 then
                     --when len/=1024DW
                        if conv_integer(tlplengthsig) /= 1 then
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                 firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                    conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                       conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                          firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                             conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                 conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + conv_integer(not((firstdwbesig(3) 
                                    xor firstdwbesig(1)) or (firstdwbesig(2) xor firstdwbesig(0)))) + 
                                       conv_integer((firstdwbesig(3) and firstdwbesig(0)) and (firstdwbesig(2) nor 
                                          firstdwbesig(1))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                             (firstdwbesig(2) nand firstdwbesig(1))) - conv_integer(firstdwbesig(3) and 
                                                firstdwbesig(2) and firstdwbesig(1) and firstdwbesig(0)), 12);
                        end if;
                     else
                     --when len=1024DW
                        if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + conv_integer(firstdwbesig(2) 
                                    or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(2) or lastdwbesig(3)) + 
                                       conv_integer(firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(1) or 
                                          lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(0) or lastdwbesig(1) or lastdwbesig(2) or 
                                                lastdwbesig(3))), 12);
                        else
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                        end if;
                     end if;
                     tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= requesteridsig;
                     tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= tagsig;
                     tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= tlptcsig;
                     tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                        blk_function_number;
                     tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpattrsig;
                     tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                     tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                     rdreq <= '1';
                     --if blk_lnk_up = '0' then
                     --   s_axis_cr_tready_sig <= '0';
                     --   rdreqsmsig  <= init;
                     --else
                     rdreqsmsig  <= memrdreq;
                     s_axis_cr_tready_sig <= '1';
                     --end if;
                     rdreqpipelineincr <= '1';
                     rdtargetpipeline <= rdtargetpipeline + 1;
                     if (orrdreqpipeline /= rdtargetpipeline) and
                     (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                        wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                     else
                        wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                     end if;
                     s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tusersigtemp;
                  end if;
               else
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
               end if;
            
            when throttle_nd =>
               -- Nam - extremely hard to hit case
               -- coverage off -item b 1 -allfalse
               if blk_lnk_up_latch = '1' then
                  if rdndreqpipeline /= "100" then
                    --pipeline full for Cpl (i.e., compl without data - no barhit or zero len)
                     --if blk_lnk_up = '0' then
                     --   s_axis_cr_tready_sig <= '0';
                     --   rdreqsmsig  <= init;
                     --else
                     rdreqsmsig  <= memrdreq;
                     s_axis_cr_tready_sig <= '1';
                     --end if;
                     if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend or 
                       badreadreq = '1' then
                        wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                     else
                        wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                     end if;
                     tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlptcsig;
                     tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlpattrsig;
                     tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= requesteridsig;
                     tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                        blk_function_number;
                     tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= tagsig;
                     rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= rdndtlpaddrlow;
                     if badreadreq = '1' then
                        cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                     elsif zerolenreadreq = '1' then
                        cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                     end if;
                     rdndtargetpipeline <= rdndtargetpipeline +1;
                     rdndreqpipelineincr <= '1';
                     badreadreq <= '0';
                     zerolenreadreq <= '0';
                     -- NAM / JRH Tool bug doesn't exclude the second condition. removed cov off item b 2. Moved cov off.
                     if conv_integer(tlplengthsig) /= 0 then
                     --when len/=1024DW
                        -- coverage off -item b 1
                        if conv_integer(tlplengthsig) /= 1 then
                           -- Not hit for EP, include for RC
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                 firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                    conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                       conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                          firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3)) + 
                                             conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or lastdwbesig(1) or 
                                                lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                 conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + conv_integer(not((firstdwbesig(3) 
                                    xor firstdwbesig(1)) or (firstdwbesig(2) xor firstdwbesig(0)))) + conv_integer((firstdwbesig(3) 
                                       and firstdwbesig(0)) and (firstdwbesig(2) nor firstdwbesig(1))) + 
                                          conv_integer((firstdwbesig(3) and firstdwbesig(0)) and (firstdwbesig(2) nand 
                                             firstdwbesig(1))) - conv_integer(firstdwbesig(3) and firstdwbesig(2) and 
                                                firstdwbesig(1) and firstdwbesig(0)), 12);
                        end if;
                     -- NAM / JRH Tool bug doesn't exclude the second condition. Moved cov off.
                     -- coverage off
                     else
                     --when len=1024DW
                           -- Not hit for EP, include for RC
                        if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or 
                                 firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + conv_integer(firstdwbesig(2) 
                                    or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(2) or lastdwbesig(3)) + 
                                       conv_integer(firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(1) or 
                                          lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + 
                                             conv_integer(lastdwbesig(0) or lastdwbesig(1) or lastdwbesig(2) or 
                                                lastdwbesig(3))), 12);
                        else
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                        end if;
                        -- coverage on
                     end if;
                  end if;
               -- Nam - extremely hard to hit case
               -- coverage off
               else
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
               end if;
               -- coverage on
               
            -- coverage off
            when others => 
               rdreqsmsig <= init;
            -- coverage on
         end case;
         if blk_lnk_up_latch = '0' and cpltargetpipeline /= ctargetpipeline then
            rdtargetpipeline <= addrstreampipeline;
         end if;
      end if;
   end if;
end process;

cplnd_master_egress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         cplndtlpsmsig <= memcplcrtdatabeat1;
         cplndtargetpipeline <= "000";
         rdndreqpipelinedecr <= '0';
         m_axis_cc_tvalid_nd <= '0';
         m_axis_cc_tdata_nd <= (others => '0');
         m_axis_cc_tstrb_nd <= (others => '0');
         m_axis_cc_tlast_nd <= '0';
         dis_valid_nd <= '0';
         orcplndpipeline <= (others => '0');
         cplndpendcpl <= (others => '0');
      else
         if orcplndpipeline /= rdndtargetpipeline then
            cplndpendcpl(conv_integer(orcplndpipeline(1 downto 0))) <= '0';
            if master_wr_idle = '1' or wrpendflush(conv_integer(orcplndpipeline(1 downto 0)))(2 downto 0) = wrreqcomp
                       or wrpendflush(conv_integer(orcplndpipeline(1 downto 0)))(3) = '1' then
               cplndpendcpl(conv_integer(orcplndpipeline(1 downto 0))) <= '1';
               orcplndpipeline <= orcplndpipeline + 1;
            end if;
         end if;
        
         -- cplndpendcpl needs to be reset on link down event
         if blk_lnk_up_latch = '0' then
            cplndpendcpl <= (others => '0');
         end if;
         case cplndtlpsmsig is
            when memcplcrtdatabeat1 =>
               rdndreqpipelinedecr <= '0';
               m_axis_cc_tvalid_nd <= '0';
               m_axis_cc_tlast_nd <= '0';
               m_axis_cc_tstrb_nd <= x"00";
               if cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline then
                  if blk_lnk_up_latch = '1' then
                     if cplndpendcpl(conv_integer(cplndtargetpipeline(1 downto 0))) = '1' then
                        if cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) = "000" then
                           m_axis_cc_tdata_nd <= tlpndcompleterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                              cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & x"001" & '0' & "10" & "01010"
                                & '0' & tlpndtc(conv_integer(cplndtargetpipeline(1 downto 0))) & "0000" & '0' & '0' & 
                                  tlpndattr(conv_integer(cplndtargetpipeline(1 downto 0))) & "00" & "0000000001";
                        -- coverage off
                        else
                           m_axis_cc_tdata_nd <= tlpndcompleterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                              cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                                 tlpndbytecount(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & "00" & "01010" & '0' 
                                    & tlpndtc(conv_integer(cplndtargetpipeline(1 downto 0))) & "0000" & '0' & '0' & 
                                       tlpndattr(conv_integer(cplndtargetpipeline(1 downto 0))) & "00" & "0000000000";
                        -- coverage on
                        end if;
                        m_axis_cc_tstrb_nd <= (others => '1');
                        m_axis_cc_tvalid_nd <= '1';
                        if m_axis_cc_tready = '1' and m_axis_cc_tvalid_nd = '1' then
                             cplndtlpsmsig <= transfer_complete;
                             m_axis_cc_tlast_nd <= '1';
                             m_axis_cc_tdata_nd <= x"00000000" & tlpndrequesterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                tlpndtag(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                                   rdndtlpaddrl(conv_integer(cplndtargetpipeline(1 downto 0)));
                             if cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) = "000" then
                                m_axis_cc_tstrb_nd <= x"FF";
                             -- coverage off
                             else
                                m_axis_cc_tstrb_nd <= x"0F";
                             -- coverage on
                             end if;
                        --else
                        --   cplndtlpsmsig <= memcplcrtdatabeat1;
                        end if;
                     end if;

                  -- Nam - extremely hard to hit case
                  -- coverage off                         
                  else
                     cplndtlpsmsig       <= memcplcrtdatabeat1;
                     rdndreqpipelinedecr <= '1';
                     cplndtargetpipeline <= cplndtargetpipeline + 1;
                  end if;
                  --coverage on
               end if;
            
            when transfer_complete =>
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tvalid_nd <= '0';
                  m_axis_cc_tlast_nd <= '0';
                  m_axis_cc_tstrb_nd <= x"00";
                  cplndtlpsmsig <= memcplcrtdatabeat1;
                  rdndreqpipelinedecr <= '1';
                  cplndtargetpipeline <= cplndtargetpipeline + 1;
               end if;
            
         -- coverage off
         when others =>
            cplndtlpsmsig <= memcplcrtdatabeat1;
         -- coverage on
      end case;
      end if;
   end if;
end process;

cpl_master_egress: process (aclk)
variable tlplengthcntr_var : std_logic_vector(9 downto 0);
begin
   if rising_edge(aclk) then
      if reset = '0' then
         cpltlpsmsig <= memcplpipeline;
         cpltargetpipeline <= (others => '0');
         rdreqpipelinedecr <= '0';
         cplpacket1 <= '0';
         m_axis_cc_tdatatemp64 <= (others=>'0');
         firstdwen   <= '0';
         lnkdowndataflush <= '0';
         m_axis_cc_tvalid_d <= '0';
         m_axis_cc_tstrb_d <= (others => '0');
         m_axis_cc_tlast_d <= '0';
         rd_en_sig <= '0';
         cplcounter <= (others => '0');
         cpldsplitcounttemp <= (others => '0');
         rdtlpaddrltemp <= (others => '0');
         ctlpbytecounttemp <= (others => '0');
         ctlplengthtemp <= (others => '0');
         tlplengthcntr <= (others => '0');
         tlplengthcntr_var := (others => '0');
         dis_valid_d <= '0';
         m_axis_cc_tdata_h <= (others => '0');
         data_phase <= '0';
         dis_rden <= '0';
         corruptdataflush <= '0';
         wait_till_not_empty <= '0';
         totallength <= (others => '0');
         totalbytecount <= (others => '0');
         linkdownflushdepth <= (others => '0');
         rrespdelayed <= '0';
      else
         case cpltlpsmsig is
            when memcplpipeline =>
               rdreqpipelinedecr <= '0';
               m_axis_cc_tlast_d <= '0';
               rd_en_sig <= '0';
               m_axis_cc_tstrb_d <= x"00";
               m_axis_cc_tvalid_d <= '0';
               if blk_lnk_up_latch = '1' then
                  if cplndtargetpipeline = rdndtargetpipeline then
                     if cpltargetpipeline /= ctargetpipeline then
                        cplcounter <= "00000";
                        cpldsplitcounttemp <= cpldsplitcount(conv_integer(cpltargetpipeline(1 downto 0)));
                        ctlpbytecounttemp <= ctlpbytecount0(conv_integer(cpltargetpipeline(1 downto 0)));
                        ctlplengthtemp <= ctlplength0(conv_integer(cpltargetpipeline(1 downto 0)));
                        totallength <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
                        tlplengthcntr_var := 
                          conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                            conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(2)))/2 + 
                              (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                                conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(2))) mod 2, 10);
                        if tlplengthcntr_var = "0000000000" then
                           linkdownflushdepth <= "1000000000";
                        else
                           linkdownflushdepth <= tlplengthcntr_var;
                        end if;
                        totalbytecount <= tlpbytecount(conv_integer(cpltargetpipeline(1 downto 0)));
                        cplpacket1 <= '1';
                        rdtlpaddrltemp <= rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)));
                        cpltlpsmsig <= memcplcrtdatabeat1;
                        rrespdelayed <= '0';
                     else
                        cpltlpsmsig <= memcplpipeline;
                     end if;
                  end if;
               -- Nam - extremely hard to hit case - we covered this in the weekend run with 10 hits
               -- coverage off                      
               elsif cpltargetpipeline /= ctargetpipeline and empty = '0' then
                  cpltlpsmsig <= blklinkdown_corruptdata;
                  lnkdowndataflush <= '1';
                  tlplengthcntr <= 
                     conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                        conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(2)))/2 + 
                           (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                              conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(2))) mod 2, 10);
                  rd_en_sig <= '1';
               end if;
               -- coverage on
            when memcplcrtdatabeat1 =>
               m_axis_cc_tlast_d <= '0';
               rd_en_sig <= '0';
               rrespdelayed <= rresp(conv_integer(cpltargetpipeline(1 downto 0)))(2);
                  if (((cplpendcpl(conv_integer(cpltargetpipeline(1 downto 0))) = '1' and rrespdelayed = '1') or 
                     slv_write_idle = '1') and rresp(conv_integer(cpltargetpipeline(1 downto 0)))(2) = '1')
                     or blk_lnk_up_latch = '0' then
                  --ordering & rresp check
                     if rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1 downto 0) = "00" then
                        if blk_lnk_up_latch = '1' then
                           m_axis_cc_tdata_h <= tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                 rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0))
                                 & '0' & (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                    rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & ctlpbytecounttemp & '0' & "10" &
                                       "01010" & '0' & tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & '0' & '0' & 
                                          tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & ctlplengthtemp;
                           tlplengthcntr <= conv_std_logic_vector((conv_integer(ctlplengthtemp))/2, 10);
                           m_axis_cc_tstrb_d <= (others => '1');
                           m_axis_cc_tvalid_d <= not(empty);
                           if (m_axis_cc_tready = '1' and m_axis_cc_tvalid_d = '1') then
                              if cplpacket1 = '0' then
                                 m_axis_cc_tdata_h <= little_to_big_endian32(dout(31 downto 0)) & 
                                    tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0)))
                                       & tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & x"00";
                              else
                                 if rdtlpaddrltemp(2) /= '1' then
                                    m_axis_cc_tdata_h <= little_to_big_endian32(dout(31 downto 0)) & 
                                       tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0)))
                                          & tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp;
                                 else
                                    m_axis_cc_tdata_h <= little_to_big_endian32(dout(63 downto 32)) & 
                                       tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0)))
                                          & tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp;
                                 end if;
                              end if;
                              m_axis_cc_tdatatemp64 <= dout(63 downto 32);
                              rd_en_sig <= '1';
                              if ctlplengthtemp = "0000000001" then
                                 m_axis_cc_tlast_d <= '1';
                                 if cplcounter = cpldsplitcounttemp then
                                 cpltlpsmsig <= memcpltxonedw;
                                 else
                                 cpltlpsmsig <= memcpltxdata;
                                 end if;
                              else
                                 cpltlpsmsig <= memcpltxdata;
                              end if;
                              linkdownflushdepth <= linkdownflushdepth - conv_std_logic_vector((conv_integer(ctlplengthtemp))/2 + 
                                conv_integer(ctlplengthtemp(0)), 10);
                           --else
                           --   cpltlpsmsig <= memcplcrtdatabeat1;
                           end if;
                        else
                           if empty = '0' then
                              cpltlpsmsig       <= blklinkdown_corruptdata;
                              m_axis_cc_tvalid_d <= '0';
                              tlplengthcntr <= linkdownflushdepth;
                              rd_en_sig            <= '1';
                              lnkdowndataflush <= '1';
                           else
                              cpltlpsmsig       <= memcplpipeline;
                           end if;
                        end if;
                     else
                        if blk_lnk_up_latch = '1' then
                           m_axis_cc_tdata_h <= tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                 rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0))
                                    & '0' & (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                       rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & totalbytecount & '0' & 
                                          "00" & "01010" & '0' & tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & 
                                             '0' & '0' & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & totallength;
                           m_axis_cc_tstrb_d <= (others => '1');
                           m_axis_cc_tvalid_d <= '1';
                           if m_axis_cc_tready = '1' and m_axis_cc_tvalid_d = '1' then
                                m_axis_cc_tdata_h <= x"00000000" & tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                   tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp;
                                cpltlpsmsig <= blklinkdown_corruptdata;
                                corruptdataflush <= '1';
                                tlplengthcntr <= 
                                   conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                                      conv_integer(rdtlpaddrltemp(2)))/2 + 
                                         (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                                            conv_integer(rdtlpaddrltemp(2))) mod 2, 10);
                                rd_en_sig <= '1';
                                m_axis_cc_tlast_d <= '1';
                                m_axis_cc_tstrb_d <= x"0F";
                           --else
                           --   cpltlpsmsig <= memcplcrtdatabeat1;
                           end if;
                           
                        -- Nam - extremely hard to hit case
                        -- coverage off                               
                        else
                           if empty = '0' then
                              cpltlpsmsig       <= blklinkdown_corruptdata;
                              m_axis_cc_tvalid_d <= '0';
                              tlplengthcntr <= 
                                 conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                                    conv_integer(rdtlpaddrltemp(2)))/2 + 
                                       (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                                          conv_integer(rdtlpaddrltemp(2))) mod 2, 10);
                              rd_en_sig            <= '1';
                              lnkdowndataflush <= '1';
                           else
                              cpltlpsmsig       <= memcplpipeline;
                           end if;
                        end if;
                        -- coverage on
                     end if;
                  end if;
            
            when blklinkdown_corruptdata =>
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tvalid_d <= '0';
               end if;
               rdreqpipelinedecr <= '0';
               if empty = '0' then
               wait_till_not_empty <= '1';
               if tlplengthcntr /= "0000000001" then
                  -- CR 653816:
                  -- 1024DW data for read request requires 200 beats to flush out data from FIFO
                  -- One beat contains two DWs so tlplengthcntr has to be adjusted to "1FF"
                  if tlplengthcntr = "0000000000" then
                     tlplengthcntr <= "0111111111";
                  else
                     tlplengthcntr <= tlplengthcntr - 1;
                  end if;
                  rd_en_sig <= '1';
               else
                  if lnkdowndataflush = '1' then
                     if cpltargetpipeline + 1 /= ctargetpipeline then
                           tlplengthcntr <= 
                           conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)+1))) + 
                              conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)+1))(2)))/2 + 
                                 (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)+1))) + 
                                    conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)+1))(2))) mod 2, 10);
                        --rdreqpipelinedecr <= '1';
                        cpltargetpipeline <= cpltargetpipeline + 1;
                     else
                        -- Nam - enhance bridge doesn't throttle
                        -- coverage off -item bc 1 -allfalse -condrow 3
                        if m_axis_cc_tvalid_d = '0' or m_axis_cc_tready = '1' then
                           cpltlpsmsig <= memcplpipeline;
                           --rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                           wait_till_not_empty <= '0';
                        end if;
                        rd_en_sig <= '0';
                        lnkdowndataflush <= '0';
                     end if;
                  else
                     -- Nam - enhance bridge doesn't throttle
                     -- coverage off -item bc 1 -allfalse -condrow 3
                     if m_axis_cc_tvalid_d = '0' or m_axis_cc_tready = '1' then
                        cpltlpsmsig <= memcplpipeline;
                        rdreqpipelinedecr <= '1';
                        cpltargetpipeline <= cpltargetpipeline + 1;
                        wait_till_not_empty <= '0';
                     end if;
                     rd_en_sig <= '0';
                     corruptdataflush <= '0';
                  end if;
               end if;
               end if;
            
            when memcpltxonedw =>
               -- Nam - enhance bridge doesn't throttle
               -- coverage off -item b 1 -allfalse            
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tvalid_d <= '0';
                  rd_en_sig <= '0';
                  m_axis_cc_tlast_d <= '0';
                  cpltlpsmsig <= memcplpipeline;
                  rdreqpipelinedecr <= '1';
                  cpltargetpipeline <= cpltargetpipeline + 1;
               end if;
            
            when memcpltxdata =>
               if empty = '0' or tlplengthcntr = "0000000000" then
                  -- Nam - enhance bridge doesn't throttle
                  -- coverage off -item b 1 -allfalse
                  if m_axis_cc_tready = '1' then
                     rd_en_sig <= '0';
                     m_axis_cc_tvalid_d <= not(empty);
                     data_phase <= '1';
                     m_axis_cc_tdatatemp64 <= dout(63 downto 32);
                     if tlplengthcntr = "0000000001" then
                        m_axis_cc_tlast_d <= '1';
                        if (conv_integer(ctlplengthtemp) + 1) mod 2 = 0 then
                           m_axis_cc_tstrb_d <= x"FF";
                        else
                           m_axis_cc_tstrb_d <= x"0F";
                           if rdtlpaddrltemp(2) = '0' or cplpacket1 = '0' then
                              dis_rden <= '1';
                           end if;
                        end if;
                     end if;
                     if tlplengthcntr = "0000000000" then
                        data_phase <= '0';
                        dis_rden <= '0';
                        m_axis_cc_tvalid_d <= '0';
                        m_axis_cc_tlast_d <= '0';
                        m_axis_cc_tstrb_d <= x"00";
                        if cplcounter /= cpldsplitcounttemp then
                           cpltlpsmsig <= memcplcrtdatabeat1;
                           cplcounter <= cplcounter + 1;
                           if cplcounter /= "00000" then
                              ctlpbytecounttemp <= ctlpbytecounttemp - 
                                 (ctlplength1(conv_integer(cpltargetpipeline(1 downto 0))) & "00");
                           else
                              ctlpbytecounttemp <= ctlpbytecounttemp - 
                                 ctlpbytecount1(conv_integer(cpltargetpipeline(1 downto 0)));
                           end if;
                           if cplcounter+1 /= cpldsplitcounttemp then
                              ctlplengthtemp <= ctlplength1(conv_integer(cpltargetpipeline(1 downto 0)));
                           else
                              ctlplengthtemp <= ctlplength2(conv_integer(cpltargetpipeline(1 downto 0)));
                           end if;
                           cplpacket1 <= '0';
                        else
                           cpltlpsmsig <= memcplpipeline;
                           rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                        end if;
                     else
                        tlplengthcntr <= tlplengthcntr - 1;
                     end if;
                  end if;
               end if;
         
            -- coverage off
            when others =>
               cpltlpsmsig <= memcplpipeline;
            -- coverage on
         end case;
         --if blk_lnk_up = '0' and blk_lnk_up_d = '1' then
         --   cpltargetpipeline <= cpltargetpipeline - rdreqpipeline;
         --end if;
      end if;
   end if;
end process;
end generate;

data_width_128: if C_S_AXIS_DATA_WIDTH = 128 generate
rd_master_ingress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cr_tready_sig    <= '0';
         rdreqpipelineincr   <= '0';
         rdtargetpipeline    <= (others => '0');
         tlplengthsig        <= (others => '0');
         firstdwbesig        <= (others => '0');
         lastdwbesig         <= (others => '0');
         tlpaddrhigh         <= (others => '0');
         tlpaddrlow          <= (others => '0');
         tlpfmtsig           <= (others => '0');
         rdreqsmsig          <= init;
         rdreq               <= '0';
         badreadreq          <= '0';
         zerolenreadreq      <= '0';
         rdndreqpipelineincr <= '0';
         rdndtargetpipeline  <= "000";
         s_axis_cr_tusersig <= (others => (others => '0'));
         s_axis_cr_tusersigtemp <= (others => '0');
      else
         case rdreqsmsig is
            when init =>
               if lnkdowndataflush = '0' and blk_lnk_up_latch = '1' then
                  s_axis_cr_tready_sig <= '1';
                  rdreqsmsig       <= memrdreq;
               end if;
            
            when memrdreq =>
               rdreqpipelineincr <= '0';
               rdndreqpipelineincr <= '0';
               rdreq <= '0';
               if blk_lnk_up_latch = '1' then
                  if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                     if s_axis_cr_tdata(30) = '0' then
                        if s_axis_cr_tdata(28 downto 24) = "00000" then
                           tlpattrsig <= s_axis_cr_tdata(13 downto 12);
                           tlplengthsig <= s_axis_cr_tdata(9 downto 0);
                           tlptcsig     <= s_axis_cr_tdata(22 downto 20);
                           lastdwbesig  <= s_axis_cr_tdata(39 downto 36);
                           firstdwbesig <= s_axis_cr_tdata(35 downto 32);
                           requesteridsig  <= s_axis_cr_tdata(63 downto 48);
                           tagsig          <= s_axis_cr_tdata(47 downto 40);
                           if s_axis_cr_tdata(29) = '0' then
                              if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                                 if ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '1') or (C_PCIEBAR_NUM > 1 and (s_axis_cr_tuser(2) = 
                                    '1' or s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) 
                                    and s_axis_cr_tdata(35 downto 32) /= "0000" then
                                    if rdreqpipeline /= "100" then
                                       tlpaddrlow <= s_axis_cr_tdata(95 downto 66) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or 
                                               s_axis_cr_tdata(32))) + conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) 
                                                 or s_axis_cr_tdata(33) or s_axis_cr_tdata(32)))), 2);
                                       tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(95 downto 66) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(95 downto 66) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(70 downto 66) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 0 then
                                          if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 1 then
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(9 downto 0)-2)*4 + 
                                                  (conv_integer(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or
                                                    s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(39)) + 
                                                      conv_integer(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or 
                                                        s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38) or 
                                                          s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                            s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                              s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                                conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36)
                                                                  or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                    s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(35)) + 
                                                  conv_integer(s_axis_cr_tdata(34)) + conv_integer(s_axis_cr_tdata(33)) + 
                                                    conv_integer(s_axis_cr_tdata(32)) + conv_integer(not((s_axis_cr_tdata(35) xor 
                                                      s_axis_cr_tdata(33)) or (s_axis_cr_tdata(34) xor s_axis_cr_tdata(32)))) + 
                                                        conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                          (s_axis_cr_tdata(34) nor s_axis_cr_tdata(33))) + 
                                                            conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                              (s_axis_cr_tdata(34) nand s_axis_cr_tdata(33))) - 
                                                                conv_integer(s_axis_cr_tdata(35) and s_axis_cr_tdata(34) and 
                                                                  s_axis_cr_tdata(33) and s_axis_cr_tdata(32)), 12);
                                          end if;
                                       else
                                          if s_axis_cr_tdata(32) /= '1' or s_axis_cr_tdata(39) /= '1' then
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(s_axis_cr_tdata(35) or 
                                                  s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32)) + 
                                                    conv_integer(s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(34) or 
                                                      s_axis_cr_tdata(33) or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38)
                                                        or s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                          s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                            s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                              conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36) 
                                                                or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                  s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                                          end if;
                                       end if;
                                       tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(63 downto 48);
                                       tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(47 downto 40);
                                       tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(22 downto 20);
                                       tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & 
                                          blk_device_number & blk_function_number;
                                       tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(13 downto 12);
                                       tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(9 downto 0);
                                       tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(9 downto 0);
                                       rdreq <= '1';
                                       rdreqsmsig  <= memrdreq;
                                       rdreqpipelineincr <= '1';
                                       rdtargetpipeline <= rdtargetpipeline + 1;
                                       if (orrdreqpipeline /= rdtargetpipeline) and
                                       (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                                          wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                                       else
                                          wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                                       end if;
                                       if C_PCIEBAR_AS = 0 then
                                          s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(C_PCIEBAR_NUM-1 downto 0) 
                                             <= s_axis_cr_tuser(C_PCIEBAR_NUM+1 downto 2);
                                       else
                                          for i in 0 to C_PCIEBAR_NUM-1 loop
                                             s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(i) <= 
                                                s_axis_cr_tuser(2*(i+1));
                                          end loop;
                                       end if;
                                    else
                                       rdreqsmsig   <= throttle;
                                       s_axis_cr_tready_sig <= '0';
                                       rdreq <= '0';
                                       tlpaddrlow <= s_axis_cr_tdata(95 downto 66) & 
                                          conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                            conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                              conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32)))
                                                + conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33)
                                                  or s_axis_cr_tdata(32)))), 2);
                                       if C_PCIEBAR_AS = 0 then
                                          s_axis_cr_tusersigtemp(C_PCIEBAR_NUM-1 downto 0) <= 
                                             s_axis_cr_tuser(C_PCIEBAR_NUM+1 downto 2);
                                       else
                                          for i in 0 to C_PCIEBAR_NUM-1 loop
                                             s_axis_cr_tusersigtemp(i) <= s_axis_cr_tuser(2*(i+1));
                                          end loop;
                                       end if;
                                    end if;
                                 else
                                    if rdndreqpipeline /= "100" then
                                       if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend
                                         or badreadreq = '1' then
                                          wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                                       else
                                          wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                                       end if;
                                       tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(22 downto 20);
                                       tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(13 downto 12);
                                       tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                          s_axis_cr_tdata(63 downto 48);
                                       tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & 
                                          blk_device_number & blk_function_number;
                                       tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(47 downto 40);
                                       rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(70 downto 66) 
                                         & conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or 
                                               s_axis_cr_tdata(32))) + conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) 
                                                 or s_axis_cr_tdata(33) or s_axis_cr_tdata(32)))), 2);
                                       if ((s_axis_cr_tuser(2) = '0' and C_PCIEBAR_NUM = 1) or (C_PCIEBAR_NUM > 1 and s_axis_cr_tuser(2) = '0' 
                                          and s_axis_cr_tuser(3) = '0' and s_axis_cr_tuser(4) = '0' and s_axis_cr_tuser(6) = '0')) then
                                          cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                                       elsif s_axis_cr_tdata(35 downto 32) = "0000" then
                                          cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                                       end if;
                                       rdndtargetpipeline <= rdndtargetpipeline +1;
                                       rdndreqpipelineincr <= '1';
                                       if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 0 then
                                          if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 1 then
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(9 downto 0)-2)*4 + 
                                                  (conv_integer(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                    or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(39)) + 
                                                      conv_integer(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or 
                                                        s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38) or 
                                                          s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                            s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                              s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                                conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36)
                                                                  or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                    s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                               conv_std_logic_vector(conv_integer(s_axis_cr_tdata(35)) + 
                                                 conv_integer(s_axis_cr_tdata(34)) + conv_integer(s_axis_cr_tdata(33)) + 
                                                   conv_integer(s_axis_cr_tdata(32)) + conv_integer(not((s_axis_cr_tdata(35) xor 
                                                     s_axis_cr_tdata(33)) or (s_axis_cr_tdata(34) xor s_axis_cr_tdata(32)))) + 
                                                       conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                         (s_axis_cr_tdata(34) nor s_axis_cr_tdata(33))) + 
                                                           conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                             (s_axis_cr_tdata(34) nand s_axis_cr_tdata(33))) - 
                                                               conv_integer(s_axis_cr_tdata(35) and s_axis_cr_tdata(34) and 
                                                                 s_axis_cr_tdata(33) and s_axis_cr_tdata(32)), 12);
                                          end if;
                                       else
                                          if s_axis_cr_tdata(32) /= '1' and s_axis_cr_tdata(39) /= '1' then
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(s_axis_cr_tdata(35) or 
                                                  s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32)) + 
                                                    conv_integer(s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(34) or 
                                                      s_axis_cr_tdata(33) or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38)
                                                        or s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                          s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                            s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                              conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36) 
                                                                or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                  s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                                          end if;
                                       end if;
                                    else
                                       s_axis_cr_tready_sig <= '0';
                                       rdreqsmsig   <= throttle_nd;
                                       if ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '0') or (C_PCIEBAR_NUM > 1 and s_axis_cr_tuser(2) = '0' 
                                          and s_axis_cr_tuser(3) = '0' and s_axis_cr_tuser(4) = '0' and s_axis_cr_tuser(6) = '0')) then
                                          badreadreq <= '1';
                                       elsif s_axis_cr_tdata(35 downto 32) = "0000" then
                                          zerolenreadreq <= '1';
                                       end if;
                                       rdndtlpaddrlow <= s_axis_cr_tdata(70 downto 66) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                    end if;
                                    rdreq <= '0';
                                 end if;
                              else
                                 rdreq <= '0';
                              end if;
                           else
                              if s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                                 if ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '1' ) or (C_PCIEBAR_NUM > 1 and (s_axis_cr_tuser(2) = '1' or
                                    s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) and 
                                    s_axis_cr_tdata(35 downto 32) /= "0000" then
                                    if rdreqpipeline /= "100" then
                                       tlpaddrlow <= s_axis_cr_tdata(127 downto 98) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(127 downto 98) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(127 downto 98) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(102 downto 98) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                          conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                            conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                              conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                or s_axis_cr_tdata(32)))), 2);
                                       if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 0 then
                                          if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 1 then
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(9 downto 0)-2)*4 + 
                                                  (conv_integer(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                    or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(39)) + 
                                                      conv_integer(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or 
                                                        s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38) or 
                                                          s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                            s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                              s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                                conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36)
                                                                  or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                    s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(35)) + 
                                                  conv_integer(s_axis_cr_tdata(34)) + conv_integer(s_axis_cr_tdata(33)) + 
                                                    conv_integer(s_axis_cr_tdata(32)) + conv_integer(not((s_axis_cr_tdata(35) xor 
                                                      s_axis_cr_tdata(33)) or (s_axis_cr_tdata(34) xor s_axis_cr_tdata(32)))) + 
                                                        conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                          (s_axis_cr_tdata(34) nor s_axis_cr_tdata(33))) + 
                                                            conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                              (s_axis_cr_tdata(34) nand s_axis_cr_tdata(33))) - 
                                                                conv_integer(s_axis_cr_tdata(35) and s_axis_cr_tdata(34) and 
                                                                  s_axis_cr_tdata(33) and s_axis_cr_tdata(32)), 12);
                                          end if;
                                       else
                                          if s_axis_cr_tdata(32) /= '1' or s_axis_cr_tdata(39) /= '1' then
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(s_axis_cr_tdata(35) or 
                                                  s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))
                                                    + conv_integer(s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(34) or 
                                                      s_axis_cr_tdata(33) or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38)
                                                        or s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                          s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                            s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                              conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36) 
                                                                or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                  s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                                          end if;
                                       end if;
                                       tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(63 downto 48);
                                       tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(47 downto 40);
                                       tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(22 downto 20);
                                       tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & 
                                          blk_device_number & blk_function_number;
                                       tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(13 downto 12);
                                       tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(9 downto 0);
                                       tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(9 downto 0);
                                       rdreq <= '1';
                                       rdreqsmsig  <= memrdreq;
                                       rdreqpipelineincr <= '1';
                                       rdtargetpipeline <= rdtargetpipeline + 1;
                                       if (orrdreqpipeline /= rdtargetpipeline) and
                                       (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                                          wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                                       else
                                          wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                                       end if;
                                       for i in 0 to C_PCIEBAR_NUM-1 loop
                                          s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0)))(i) <= 
                                             s_axis_cr_tuser(2*(i+1));
                                       end loop;
                                    else
                                       rdreqsmsig   <= throttle;
                                       s_axis_cr_tready_sig <= '0';
                                       rdreq <= '0';
                                       tlpaddrlow <= s_axis_cr_tdata(127 downto 98) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                               or s_axis_cr_tdata(32)))), 2);
                                       for i in 0 to C_PCIEBAR_NUM-1 loop
                                          s_axis_cr_tusersigtemp(i) <= s_axis_cr_tuser(2*(i+1));
                                       end loop;
                                    end if;
                                 else
                                    if rdndreqpipeline /= "100" then
                                       rdreqsmsig  <= memrdreq;
                                       if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend
                                         or badreadreq = '1' then
                                          wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                                       else
                                          wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                                       end if;
                                       tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(22 downto 20);
                                       tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(13 downto 12);
                                       tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                          s_axis_cr_tdata(63 downto 48);
                                       tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & 
                                          blk_device_number & blk_function_number;
                                       tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(47 downto 40);
                                       rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= s_axis_cr_tdata(102 downto 98) 
                                         & conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                       if ((s_axis_cr_tuser(2) = '0' and C_PCIEBAR_NUM = 1) or (C_PCIEBAR_NUM > 1 and s_axis_cr_tuser(2) = '0'
                                          and s_axis_cr_tuser(3) = '0' and s_axis_cr_tuser(4) = '0' and s_axis_cr_tuser(6) = '0')) then
                                          cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                                       elsif s_axis_cr_tdata(35 downto 32) = "0000" then
                                          cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                                       end if;
                                       rdndtargetpipeline <= rdndtargetpipeline +1;
                                       rdndreqpipelineincr <= '1';
                                       if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 0 then
                                          if conv_integer(s_axis_cr_tdata(9 downto 0)) /= 1 then
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(9 downto 0)-2)*4 + 
                                                  (conv_integer(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                    or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(39)) + 
                                                      conv_integer(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or 
                                                        s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38) or 
                                                          s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                            s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                              s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                                conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36)
                                                                  or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                    s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(s_axis_cr_tdata(35)) + 
                                                  conv_integer(s_axis_cr_tdata(34)) + conv_integer(s_axis_cr_tdata(33)) + 
                                                    conv_integer(s_axis_cr_tdata(32)) + conv_integer(not((s_axis_cr_tdata(35) 
                                                      xor s_axis_cr_tdata(33)) or (s_axis_cr_tdata(34) xor s_axis_cr_tdata(32)))) + 
                                                        conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                          (s_axis_cr_tdata(34) nor s_axis_cr_tdata(33))) + 
                                                            conv_integer((s_axis_cr_tdata(35) and s_axis_cr_tdata(32)) and 
                                                              (s_axis_cr_tdata(34) nand s_axis_cr_tdata(33))) - 
                                                                conv_integer(s_axis_cr_tdata(35) and s_axis_cr_tdata(34) and 
                                                                  s_axis_cr_tdata(33) and s_axis_cr_tdata(32)), 12);
                                          end if;
                                       else
                                          if s_axis_cr_tdata(32) /= '1' and s_axis_cr_tdata(39) /= '1' then
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                                                conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(s_axis_cr_tdata(35) or 
                                                  s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))
                                                    + conv_integer(s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(34) or 
                                                      s_axis_cr_tdata(33) or s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(38)
                                                        or s_axis_cr_tdata(39)) + conv_integer(s_axis_cr_tdata(33) or 
                                                          s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(37) or 
                                                            s_axis_cr_tdata(38) or s_axis_cr_tdata(39)) + 
                                                              conv_integer(s_axis_cr_tdata(32)) + conv_integer(s_axis_cr_tdata(36) 
                                                                or s_axis_cr_tdata(37) or s_axis_cr_tdata(38) or 
                                                                  s_axis_cr_tdata(39))), 12);
                                          else
                                             tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                                          end if;
                                       end if;
                                    else
                                       s_axis_cr_tready_sig <= '0';
                                       rdreqsmsig   <= throttle_nd;
                                       if ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '0') or (C_PCIEBAR_NUM > 1 and s_axis_cr_tuser(2) = '0'
                                          and s_axis_cr_tuser(3) = '0' and s_axis_cr_tuser(4) = '0' and s_axis_cr_tuser(6) = '0')) then
                                          badreadreq <= '1';
                                       elsif s_axis_cr_tdata(35 downto 32) = "0000" then
                                          zerolenreadreq <= '1';
                                       end if;
                                       rdndtlpaddrlow <= s_axis_cr_tdata(102 downto 98) & 
                                         conv_std_logic_vector((conv_integer(not(s_axis_cr_tdata(32))) + 
                                           conv_integer(not(s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                             conv_integer(not(s_axis_cr_tdata(34) or s_axis_cr_tdata(33) or s_axis_cr_tdata(32))) + 
                                               conv_integer(not(s_axis_cr_tdata(35) or s_axis_cr_tdata(34) or s_axis_cr_tdata(33) 
                                                 or s_axis_cr_tdata(32)))), 2);
                                    end if;
                                    rdreq <= '0';
                                 end if;
                              else
                                 rdreq <= '0';
                              end if;
                           end if;
                        --else
                        --   rdreq <= '0';
                        end if;
                     --else
                     --   rdreq <= '0';
                     end if;
                  else
                     rdreq <= '0';
                  end if;
               elsif s_axis_cr_tvalid = '1' and s_axis_cr_tlast = '1' then
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
                  rdreq <= '0';
               end if;

            when throttle =>
               if blk_lnk_up_latch = '1' then
                  if rdreqpipeline /= "101" then
                    --pipeline full for CplD (i.e., compl with data)
                     tlpaddrl(conv_integer(rdtargetpipeline(1 downto 0)))    <= tlpaddrlow;
                     tlpaddrl_out(conv_integer(rdtargetpipeline(1 downto 0)))    <= tlpaddrlow;
                     rdtlpaddrl(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpaddrlow(6 downto 0);
                     if conv_integer(tlplengthsig) /= 0 then
                     --when len/=1024DW
                        if conv_integer(tlplengthsig) /= 1 then
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                  conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                    conv_integer(lastdwbesig(2) or lastdwbesig(3)) + 
                                      conv_integer(firstdwbesig(1) or firstdwbesig(0)) + 
                                        conv_integer(lastdwbesig(1) or lastdwbesig(2) 
                                          or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or 
                                        lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                  conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                    firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                      (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) 
                                        and (firstdwbesig(2) nand firstdwbesig(1))) - conv_integer(firstdwbesig(3) and 
                                        firstdwbesig(2) and firstdwbesig(1) and firstdwbesig(0)), 12);
                        end if;
                     else
                     --when len=1024DW
                        if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or 
                                firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + conv_integer(firstdwbesig(2) 
                                  or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(2) or lastdwbesig(3)) + 
                                    conv_integer(firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(1) or 
                                      lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + 
                                        conv_integer(lastdwbesig(0) or lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpbytecount(conv_integer(rdtargetpipeline(1 downto 0))) <= (others => '0');
                        end if;
                     end if;
                     tlprequesterid(conv_integer(rdtargetpipeline(1 downto 0))) <= requesteridsig;
                     tlptag(conv_integer(rdtargetpipeline(1 downto 0))) <= tagsig;
                     tlptc(conv_integer(rdtargetpipeline(1 downto 0))) <= tlptcsig;
                     tlpcompleterid(conv_integer(rdtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                        blk_function_number;
                     tlpattr(conv_integer(rdtargetpipeline(1 downto 0))) <= tlpattrsig;
                     tlplength(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                     tlplength_out(conv_integer(rdtargetpipeline(1 downto 0))) <= tlplengthsig;
                     --if blk_lnk_up = '0' then
                     --   s_axis_cr_tready_sig <= '0';
                     --else
                     s_axis_cr_tready_sig <= '1';
                     --end if;
                     rdreq <= '1';
                     rdreqsmsig  <= memrdreq;
                     rdreqpipelineincr <= '1';
                     rdtargetpipeline <= rdtargetpipeline + 1;
                     if (orrdreqpipeline /= rdtargetpipeline) and
                     (wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend) then
                        wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                     else
                        wrpendingsig(conv_integer(rdtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                     end if;
                     s_axis_cr_tusersig(conv_integer(rdtargetpipeline(1 downto 0))) <= s_axis_cr_tusersigtemp;
                  end if;
               else
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
               end if;
            
            when throttle_nd =>
               if blk_lnk_up_latch = '1' then
                  if rdndreqpipeline /= "101" then
                    --pipeline full for Cpl (i.e., compl without data - no barhit or zero len)
                     rdreqsmsig  <= memrdreq;
                     if wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0) - "01"))(2 downto 0) = wrreqpend
                       or badreadreq = '1' then
                        wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '1' & wrreqpend;
                     else
                        wrpendflush(conv_integer(rdndtargetpipeline(1 downto 0))) <= '0' & wrreqpend;
                     end if;
                     tlpndtc(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlptcsig;
                     tlpndattr(conv_integer(rdndtargetpipeline(1 downto 0))) <= tlpattrsig;
                     tlpndrequesterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= requesteridsig;
                     tlpndcompleterid(conv_integer(rdndtargetpipeline(1 downto 0))) <= blk_bus_number & blk_device_number & 
                        blk_function_number;
                     tlpndtag(conv_integer(rdndtargetpipeline(1 downto 0))) <= tagsig;
                     rdndtlpaddrl(conv_integer(rdndtargetpipeline(1 downto 0))) <= rdndtlpaddrlow;
                     if badreadreq = '1' then
                        cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "001";
                     elsif zerolenreadreq = '1' then
                        cplndstatuscode(conv_integer(rdndtargetpipeline(1 downto 0))) <= "000";
                     end if;
                     rdndtargetpipeline <= rdndtargetpipeline +1;
                     rdndreqpipelineincr <= '1';
                     badreadreq <= '0';
                     zerolenreadreq <= '0';
                     --if blk_lnk_up = '0' then
                     --   s_axis_cr_tready_sig <= '0';
                     --else
                     s_axis_cr_tready_sig <= '1';
                     --end if;
                     if conv_integer(tlplengthsig) /= 0 then
                     --when len/=1024DW
                        if conv_integer(tlplengthsig) /= 1 then
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(tlplengthsig-2)*4 + (conv_integer(firstdwbesig(3) or 
                                firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                  conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                    conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                      firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) 
                                        or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or 
                                          lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(firstdwbesig(3)) + conv_integer(firstdwbesig(2)) + 
                                conv_integer(firstdwbesig(1)) + conv_integer(firstdwbesig(0)) + 
                                  conv_integer(not((firstdwbesig(3) xor firstdwbesig(1)) or (firstdwbesig(2) xor 
                                    firstdwbesig(0)))) + conv_integer((firstdwbesig(3) and firstdwbesig(0)) and 
                                      (firstdwbesig(2) nor firstdwbesig(1))) + conv_integer((firstdwbesig(3) and 
                                        firstdwbesig(0)) and (firstdwbesig(2) nand firstdwbesig(1))) - 
                                          conv_integer(firstdwbesig(3) and firstdwbesig(2) and firstdwbesig(1) and 
                                            firstdwbesig(0)), 12);
                        end if;
                     else
                     --when len=1024DW
                        if firstdwbesig(0) /= '1' or lastdwbesig(3) /= '1' then
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= 
                              conv_std_logic_vector(conv_integer(1022)*4 + (conv_integer(firstdwbesig(3) or firstdwbesig(2) or 
                                firstdwbesig(1) or firstdwbesig(0)) + conv_integer(lastdwbesig(3)) + 
                                  conv_integer(firstdwbesig(2) or firstdwbesig(1) or firstdwbesig(0)) + 
                                    conv_integer(lastdwbesig(2) or lastdwbesig(3)) + conv_integer(firstdwbesig(1) or 
                                      firstdwbesig(0)) + conv_integer(lastdwbesig(1) or lastdwbesig(2) 
                                        or lastdwbesig(3)) + conv_integer(firstdwbesig(0)) + conv_integer(lastdwbesig(0) or 
                                          lastdwbesig(1) or lastdwbesig(2) or lastdwbesig(3))), 12);
                        else
                           tlpndbytecount(conv_integer(rdndtargetpipeline(1 downto 0))) <= (others => '0');
                        end if;
                     end if;
                  end if;
               else
                  rdreqsmsig       <= init;
                  s_axis_cr_tready_sig <= '0';
               end if;

            -- coverage off
            when others => 
               rdreqsmsig <= init;
            -- coverage on
         end case;
         if blk_lnk_up_latch = '0' and cpltargetpipeline /= ctargetpipeline then
            rdtargetpipeline <= addrstreampipeline;
         end if;
      end if;
   end if;
end process;

cplnd_master_egress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         cplndtlpsmsig <= memcplcrtdatabeat1;
         cplndtargetpipeline <= "000";
         rdndreqpipelinedecr <= '0';
         m_axis_cc_tvalid_nd <= '0';
         m_axis_cc_tdata_nd <= (others => '0');
         m_axis_cc_tstrb_nd <= (others => '0');
         m_axis_cc_tlast_nd <= '0';
         dis_valid_nd <= '0';
         orcplndpipeline <= (others => '0');
         cplndpendcpl <= (others => '0');
      else
         if orcplndpipeline /= rdndtargetpipeline then
            cplndpendcpl(conv_integer(orcplndpipeline(1 downto 0))) <= '0';
            if master_wr_idle = '1' or wrpendflush(conv_integer(orcplndpipeline(1 downto 0)))(2 downto 0) = wrreqcomp
                       or wrpendflush(conv_integer(orcplndpipeline(1 downto 0)))(3) = '1' then
               cplndpendcpl(conv_integer(orcplndpipeline(1 downto 0))) <= '1';
               orcplndpipeline <= orcplndpipeline + 1;
            end if;
         end if;
        
         -- cplndpendcpl needs to be reset on link down event
         if blk_lnk_up_latch = '0' then
            cplndpendcpl <= (others => '0');
         end if;
         case cplndtlpsmsig is
            when memcplcrtdatabeat1 =>
               rdndreqpipelinedecr <= '0';
               m_axis_cc_tvalid_nd <= '0';
               m_axis_cc_tlast_nd <= '0';
               m_axis_cc_tstrb_nd <= x"0000";
               if cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline then
                  if blk_lnk_up_latch = '1' then
                     if cplndpendcpl(conv_integer(cplndtargetpipeline(1 downto 0))) = '1' then
                        if cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) = "000" then
                           m_axis_cc_tdata_nd <= x"00000000" & tlpndrequesterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                              tlpndtag(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                                 rdndtlpaddrl(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                    tlpndcompleterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                       cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & x"001" & '0' & "10" & 
                                          "01010" & '0' & tlpndtc(conv_integer(cplndtargetpipeline(1 downto 0))) & "0000" & '0' & 
                                            '0' & tlpndattr(conv_integer(cplndtargetpipeline(1 downto 0))) & "00" & "0000000001";
                           m_axis_cc_tstrb_nd <= x"FFFF";
                        -- coverage off
                        else
                           m_axis_cc_tdata_nd <= x"00000000" & tlpndrequesterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                              tlpndtag(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                                rdndtlpaddrl(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                  tlpndcompleterid(conv_integer(cplndtargetpipeline(1 downto 0))) & 
                                    cplndstatuscode(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & 
                                      tlpndbytecount(conv_integer(cplndtargetpipeline(1 downto 0))) & '0' & "00" & 
                                        "01010" & '0' & tlpndtc(conv_integer(cplndtargetpipeline(1 downto 0))) & "0000" & '0' & 
                                          '0' & tlpndattr(conv_integer(cplndtargetpipeline(1 downto 0))) & "00" & "0000000000";
                           m_axis_cc_tstrb_nd <= x"0FFF";
                        -- coverage on
                        end if;
                        m_axis_cc_tvalid_nd <= '1';
                        m_axis_cc_tlast_nd <= '1';
                        if m_axis_cc_tready = '1' and m_axis_cc_tvalid_nd = '1' then
                           rdndreqpipelinedecr <= '1';
                           cplndtargetpipeline <= cplndtargetpipeline + 1;
                           
                           m_axis_cc_tvalid_nd <= '0';
                           m_axis_cc_tlast_nd <= '0';
                           m_axis_cc_tstrb_nd <= x"0000";
                        end if;
                     end if;
                  else
                     rdndreqpipelinedecr <= '1';
                     cplndtargetpipeline <= cplndtargetpipeline + 1;
                  end if;
               end if;
            
         -- coverage off
         when others =>
            cplndtlpsmsig <= memcplcrtdatabeat1;
         -- coverage on
      end case;
      end if;
   end if;
end process;

tlplength_array_val <= conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0))));
rdtlpaddrl_array_val <= conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2));
rdtlpaddrltemp_array_val <= conv_integer(rdtlpaddrltemp(3 downto 2));

tlplengthcntr_var_inst : array_arith
            port map 
            (
            din0 => tlplength_array_val,
            din1 => rdtlpaddrl_array_val,
            dout => tlplengthcntr_var_tmp
            );

tlplengthcntr_inst : array_arith
            port map 
            (
            din0 => tlplength_array_val,
            din1 => rdtlpaddrltemp_array_val,
            dout => tlplengthcntr_tmp
            );


cpl_master_egress: process (aclk)
   variable tlplengthcntr_var : std_logic_vector(9 downto 0);
begin
   if rising_edge(aclk) then
      if reset = '0' then
         cpltlpsmsig <= memcplpipeline;
         cpltargetpipeline <= (others => '0');
         rdreqpipelinedecr <= '0';
         cplpacket1 <= '0';
         m_axis_cc_tdatatemp128 <= (others=>'0');
         firstdwen   <= '0';
         lnkdowndataflush <= '0';
         m_axis_cc_tvalid_d <= '0';
         m_axis_cc_tstrb_d <= (others => '0');
         m_axis_cc_tlast_d <= '0';
         rd_en_sig <= '0';
         cplcounter <= (others => '0');
         cpldsplitcounttemp <= (others => '0');
         rdtlpaddrltemp <= (others => '0');
         ctlpbytecounttemp <= (others => '0');
         ctlplengthtemp <= (others => '0');
         tlplengthcntr <= (others => '0');
         tlplengthcntr_var := (others => '0');
         dis_valid_d <= '0';
         m_axis_cc_tdata_h <= (others => '0');
         data_phase <= '0';
         dis_rden <= '0';
         corruptdataflush <= '0';
         wait_till_not_empty <= '0';
         totallength <= (others => '0');
         totalbytecount <= (others => '0');
         linkdownflushdepth <= (others => '0');
         rrespdelayed <= '0';
      else
         case cpltlpsmsig is
            when memcplpipeline =>
               rdreqpipelinedecr <= '0';
               m_axis_cc_tlast_d <= '0';
               m_axis_cc_tstrb_d <= x"0000";
               m_axis_cc_tvalid_d <= '0';
               if blk_lnk_up_latch = '1' then
                  if cplndtargetpipeline = rdndtargetpipeline then
                     if cpltargetpipeline /= ctargetpipeline then
                        rd_en_sig <= '0';
                        cplcounter <= "00000";
                        cpldsplitcounttemp <= cpldsplitcount(conv_integer(cpltargetpipeline(1 downto 0)));
                        totallength <= tlplength(conv_integer(cpltargetpipeline(1 downto 0)));
			-- Chaitanya - Updated to help meet timing
                        --if ((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                        --  conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2))) mod 4 = 0) then
                        --   tlplengthcntr_var := 
                        --   conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                        --     conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2)))/4, 10);
                        --else
                        --   tlplengthcntr_var := 
                        --      conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                        --        conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2)))/4 
                        --         + 1, 10);
                        --end if;
                        
                        --tlplengthcntr_var := conv_std_logic_vector(chaitanya3 + chaitanya2_sel, 10);
                        tlplengthcntr_var := tlplengthcntr_var_tmp;
                        if tlplengthcntr_var = "0000000000" then
                           linkdownflushdepth <= "0100000000";
                        else
                           linkdownflushdepth <= tlplengthcntr_var;
                        end if;
                        totalbytecount <= tlpbytecount(conv_integer(cpltargetpipeline(1 downto 0)));
                        cplpacket1 <= '1';
                        rdtlpaddrltemp <= rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)));
                        ctlpbytecounttemp <= ctlpbytecount0(conv_integer(cpltargetpipeline(1 downto 0)));
                        ctlplengthtemp <= ctlplength0(conv_integer(cpltargetpipeline(1 downto 0)));
                        cpltlpsmsig <= memcplcrtdatabeat1;
                        rrespdelayed <= '0';
                     else
                        cpltlpsmsig <= memcplpipeline;
                     end if;
                  end if;
               elsif cpltargetpipeline /= ctargetpipeline and empty = '0' then
                  cpltlpsmsig <= blklinkdown_corruptdata;
                  lnkdowndataflush <= '1';
		  -- Chaitanya - Updated to help meet timing
                  --if (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                  --  conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2))) mod 4 = 0 then
                  --   tlplengthcntr <= conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                  --     conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2)))/4, 10);
                  --else
                  --   tlplengthcntr <= conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                  --     conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)))(3 downto 2)))/4 + 1, 10);
                  --end if;
                  tlplengthcntr <= tlplengthcntr_var_tmp; 
                  rd_en_sig <= '1';
               end if;
            
            when memcplcrtdatabeat1 =>
               m_axis_cc_tlast_d <= '0';
               rrespdelayed <= rresp(conv_integer(cpltargetpipeline(1 downto 0)))(2);
                  if (((cplpendcpl(conv_integer(cpltargetpipeline(1 downto 0))) = '1' and rrespdelayed = '1') or 
                    slv_write_idle = '1') and rresp(conv_integer(cpltargetpipeline(1 downto 0)))(2) = '1')
                    or blk_lnk_up_latch = '0' then
                  --ordering & rresp check
                     if rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1 downto 0) = "00" then
                        if blk_lnk_up_latch = '1' then
                           if empty = '0' then
                              if cplpacket1 <= '0' then
                                 m_axis_cc_tdata_h <= 
                                    little_to_big_endian32(dout(31 downto 0)) & 
                                      tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                       tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & x"00" & 
                                          tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                             (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                                rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                   (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                                      rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                         ctlpbytecounttemp & '0' & "10" & "01010" & '0' & 
                                                            tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & '0' & '0'
                                                               & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & 
                                                       ctlplengthtemp;
                              else
                                 if rdtlpaddrltemp(3 downto 2) = "11" then
                                    m_axis_cc_tdata_h <= 
                                    little_to_big_endian32(dout(127 downto 96)) & 
                                      tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                       tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp & 
                                          tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                             (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                                rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                   (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                                      rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                       ctlpbytecounttemp & '0' & "10" & "01010" & '0' & 
                                                          tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & '0' & '0' 
                                                             & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & 
                                                                ctlplengthtemp;
                                 elsif rdtlpaddrltemp(3) = '1' then
                                    m_axis_cc_tdata_h <= 
                                    little_to_big_endian32(dout(95 downto 64)) & 
                                      tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                       tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp & 
                                          tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                             (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                                rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                   (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                                      rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                       ctlpbytecounttemp & '0' & "10" & "01010" & '0' & 
                                                          tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & '0' & '0' 
                                                             & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & 
                                                                ctlplengthtemp;
                                 elsif rdtlpaddrltemp(2) = '1' then
                                    m_axis_cc_tdata_h <= 
                                    little_to_big_endian32(dout(63 downto 32)) & 
                                      tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                       tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp & 
                                          tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                             (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                                rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                   (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                                      rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                       ctlpbytecounttemp & '0' & "10" & "01010" & '0' & 
                                                          tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & '0' & '0' 
                                                             & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & 
                                                                ctlplengthtemp;
                                 else
                                    m_axis_cc_tdata_h <= 
                                    little_to_big_endian32(dout(31 downto 0)) & 
                                      tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                       tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp & 
                                          tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                             (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                                rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                   (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                                      rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                                       ctlpbytecounttemp & '0' & "10" & "01010" & '0' & 
                                                          tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & "0000" & '0' & '0' 
                                                             & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00" & 
                                                                ctlplengthtemp;
                                 end if;
                              end if;
                              m_axis_cc_tstrb_d <= x"FFFF";
                              m_axis_cc_tdatatemp128 <= dout(127 downto 32);
                              m_axis_cc_tvalid_d <= '1';
                              if ctlplengthtemp = "0000000001" then
                                 m_axis_cc_tlast_d <= '1';
                              end if;
                              if m_axis_cc_tready = '1' and m_axis_cc_tvalid_d = '1' then
                                 if (conv_integer(ctlplengthtemp) + 3) mod 4 = 0 then
                                    tlplengthcntr <= conv_std_logic_vector(((conv_integer(ctlplengthtemp) + 3)/4)-1, 10);
                                    linkdownflushdepth <= linkdownflushdepth - 
                                      conv_std_logic_vector(((conv_integer(ctlplengthtemp) + 3)/4), 10);
                                 else
                                    tlplengthcntr <= conv_std_logic_vector((conv_integer(ctlplengthtemp) + 3)/4, 10);
                                    linkdownflushdepth <= linkdownflushdepth - 
                                      conv_std_logic_vector(((conv_integer(ctlplengthtemp) + 3)/4), 10);
                                 end if;
                                 rd_en_sig <= '1';
                                 m_axis_cc_tvalid_d <= '0';
                                 if ctlplengthtemp = "0000000001" then
                                    if cplcounter = cpldsplitcounttemp then
                                    cpltlpsmsig <= memcpltxonedw;
                                    else
                                    cpltlpsmsig <= memcpltxdata;
                                    end if;
                                    m_axis_cc_tlast_d <= '0';
                                 else
                                    cpltlpsmsig <= memcpltxdata;
                                 end if;
                              end if;
                           end if;
                        else
                           cpltlpsmsig       <= blklinkdown_corruptdata;
                           m_axis_cc_tvalid_d <= '0';
                           tlplengthcntr <= linkdownflushdepth;
                           rd_en_sig        <= '1';
                           lnkdowndataflush <= '1';
                        end if;
                     else
                        if blk_lnk_up_latch = '1' then
                           m_axis_cc_tdata_h <= x"00000000" & tlprequesterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                              tlptag(conv_integer(cpltargetpipeline(1 downto 0))) & '0' & rdtlpaddrltemp & 
                                 tlpcompleterid(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                    (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) xor 
                                       rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & 
                                          (rresp(conv_integer(cpltargetpipeline(1 downto 0)))(1) and 
                                             rresp(conv_integer(cpltargetpipeline(1 downto 0)))(0)) & '0' & totalbytecount & '0' 
                                               & "00" & "01010" & '0' & tlptc(conv_integer(cpltargetpipeline(1 downto 0))) & 
                                                 "0000" & '0' & '0' & tlpattr(conv_integer(cpltargetpipeline(1 downto 0))) & "00"
                                                   & totallength;
                           m_axis_cc_tstrb_d <= x"0FFF";
                           m_axis_cc_tvalid_d <= '1';
                           m_axis_cc_tlast_d <= '1';
                           if m_axis_cc_tready = '1' and m_axis_cc_tvalid_d = '1' then
                              cpltlpsmsig <= blklinkdown_corruptdata;
                              corruptdataflush <= '1';
                              m_axis_cc_tvalid_d <= '0';
			      -- Chaitanya - Updated to help meet timing
                              --if (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                              --  conv_integer(rdtlpaddrltemp(3 downto 2))) mod 4 = 0 then
                              --   tlplengthcntr <= 
                              --   conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                              --     conv_integer(rdtlpaddrltemp(3 downto 2)))/4, 10);
                              --else
                              --   tlplengthcntr <= 
                              --      conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                              --        conv_integer(rdtlpaddrltemp(3 downto 2)))/4 
                              --         + 1, 10);
                              --end if;
                              tlplengthcntr <= tlplengthcntr_tmp; 
                              rd_en_sig <= '1';
                           --else
                           --   cpltlpsmsig <= memcplcrtdatabeat1;
                           end if;
                        else
                           cpltlpsmsig       <= blklinkdown_corruptdata;
                           m_axis_cc_tvalid_d <= '0';
			   -- Chaitanya - Updated to help meet timing
                           --if (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                           --  conv_integer(rdtlpaddrltemp(3 downto 2))) mod 4 = 0 then
                           --   tlplengthcntr <= 
                           --   conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                           --      conv_integer(rdtlpaddrltemp(3 downto 2)))/4, 10);
                           --else
                           --   tlplengthcntr <= 
                           --      conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)))) + 
                           --        conv_integer(rdtlpaddrltemp(3 downto 2)))/4 
                           --         + 1, 10);
                           --end if;
                           tlplengthcntr <= tlplengthcntr_tmp; 
                           rd_en_sig <= '1';
                           lnkdowndataflush <= '1';
                        end if;
                     end if;
                  end if;

            when blklinkdown_corruptdata =>
               if m_axis_cc_tready = '1' then
                  m_axis_cc_tvalid_d <= '0';
               end if;
               rdreqpipelinedecr <= '0';
               if empty = '0' then
                  wait_till_not_empty <= '1';
                  if tlplengthcntr /= "0000000001" then
                    -- CR 653816:
                    -- 1024DW data for read request requires 100 beats to flush out data from FIFO
                    -- One beat contains two DWs so tlplengthcntr has to be adjusted to "FF"
                     if tlplengthcntr = "0000000000" then
                        tlplengthcntr <= "0011111111";
                     else
                        tlplengthcntr <= tlplengthcntr - 1;
                     end if;
                     rd_en_sig <= '1';
                  else
                     if lnkdowndataflush = '1' then
                        if cpltargetpipeline + 1 /= ctargetpipeline then
			   -- Chaitanya - Updated to help meet timing
                           --if (conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)+1))) + 
                           --  conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)+1))(3 downto 2))) mod 4 = 0 then
                           --   tlplengthcntr <= 
                           --   conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)+1))) + 
                           --     conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)+1))(3 downto 2)))/4, 10);
                           --else
                           --   tlplengthcntr <= 
                           --      conv_std_logic_vector((conv_integer(tlplength(conv_integer(cpltargetpipeline(1 downto 0)+1))) + 
                           --        conv_integer(rdtlpaddrl(conv_integer(cpltargetpipeline(1 downto 0)+1))(3 downto 2)))/4 
                           --         + 1, 10);
                           --end if;
                           tlplengthcntr <= tlplengthcntr_var_tmp;
                           --rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                        else
                           if m_axis_cc_tvalid_d = '0' or m_axis_cc_tready = '1' then
                              cpltlpsmsig <= memcplpipeline;
                              --rdreqpipelinedecr <= '1';
                              cpltargetpipeline <= cpltargetpipeline + 1;
                              wait_till_not_empty <= '0';
                           end if;
                           rd_en_sig <= '0';
                           lnkdowndataflush <= '0';
                        end if;
                     else
                        if m_axis_cc_tvalid_d = '0' or m_axis_cc_tready = '1' then
                           cpltlpsmsig <= memcplpipeline;
                           rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                           wait_till_not_empty <= '0';
                        end if;
                        rd_en_sig <= '0';
                        corruptdataflush <= '0';
                     end if;
                  end if;
               end if;

            when memcpltxonedw =>
               -- Don't wait for tready to come here as transfer is already complete
               --if m_axis_cc_tready = '1' then
                  rd_en_sig <= '0';
                  cpltlpsmsig <= memcplpipeline;
                  rdreqpipelinedecr <= '1';
                  cpltargetpipeline <= cpltargetpipeline + 1;
               --end if;
            
            when memcpltxdata =>
               if empty = '0' or tlplengthcntr = "0000000000" then
                  if m_axis_cc_tready = '1' or (m_axis_cc_tready = '0' and ctlplengthtemp = "0000000001") then
                     rd_en_sig <= '0';
                     m_axis_cc_tvalid_d <= not(empty);
                     data_phase <= '1';
                     m_axis_cc_tdatatemp128 <= dout(127 downto 32);
                     if tlplengthcntr = "0000000001" then
                        m_axis_cc_tlast_d <= '1';
                           case 
                           ((conv_integer(ctlplengthtemp) + 3) mod 4) is
                           when 0 =>
                              m_axis_cc_tstrb_d <= x"FFFF";
                           when 1 =>
                              m_axis_cc_tstrb_d <= x"000F";
                              if rdtlpaddrltemp(3 downto 2) /= "11" or cplpacket1 = '0' then
                                 dis_rden <= '1';
                              end if;
                           when 2 =>
                              m_axis_cc_tstrb_d <= x"00FF"; 
                              if rdtlpaddrltemp(3 downto 2) = "01" or rdtlpaddrltemp(3 downto 2) = "00" or cplpacket1 = '0' then
                                 dis_rden <= '1';
                              end if;
                           when 3 =>
                              m_axis_cc_tstrb_d <= x"0FFF"; 
                              if rdtlpaddrltemp(3 downto 2) = "00" or cplpacket1 = '0' then
                                 dis_rden <= '1';
                              end if;
                           -- coverage off
                           when others =>
                           -- coverage on
                           end case;
                     end if;
                     if tlplengthcntr = "0000000000" then
                        dis_rden <= '0';
                        data_phase <= '0';
                        m_axis_cc_tvalid_d <= '0';
                        m_axis_cc_tlast_d <= '0';
                        if cplcounter /= cpldsplitcounttemp then
                           cpltlpsmsig <= memcplcrtdatabeat1;
                           cplcounter <= cplcounter + 1;
                           if cplcounter /= "00000" then
                              ctlpbytecounttemp <= ctlpbytecounttemp - 
                                 (ctlplength1(conv_integer(cpltargetpipeline(1 downto 0))) & "00");
                           else
                              ctlpbytecounttemp <= ctlpbytecounttemp - 
                                 ctlpbytecount1(conv_integer(cpltargetpipeline(1 downto 0)));
                           end if;
                           if cplcounter+1 /= cpldsplitcounttemp then
                              ctlplengthtemp <= ctlplength1(conv_integer(cpltargetpipeline(1 downto 0)));
                           else
                              ctlplengthtemp <= ctlplength2(conv_integer(cpltargetpipeline(1 downto 0)));
                           end if;
                           cplpacket1 <= '0';
                        else
                           cpltlpsmsig <= memcplpipeline;
                           rdreqpipelinedecr <= '1';
                           cpltargetpipeline <= cpltargetpipeline + 1;
                        end if;
                     else
                        tlplengthcntr <= tlplengthcntr - 1;
                     end if;
                  end if;
               end if;
         
         -- coverage off
         when others =>
            cpltlpsmsig <= memcplpipeline;
         -- coverage on
      end case;
      end if;
   end if;
end process;
end generate;

rd_req_32_64: if C_S_AXIS_DATA_WIDTH /= 128 generate
rd_req_pipeline: process(aclk)
begin
   --pipeline buffer availability up/counter counter - CplD
   if rising_edge(aclk) then
      if reset = '0' or blk_lnk_up = '0' then
      --if reset = '0' then
         rdreqpipeline <= (others => '0');
      elsif rdreqpipelineincr = '1' and rdreqpipelinedecr = '1' then
         rdreqpipeline <= rdreqpipeline;
      elsif rdreqpipelineincr = '1' then
         rdreqpipeline <= rdreqpipeline + 1;
      elsif rdreqpipelinedecr = '1' then
         rdreqpipeline <= rdreqpipeline - 1;
      end if;
   end if;
   --pipeline buffer availability up/counter counter - Cpl
   if rising_edge(aclk) then
      if reset = '0' or blk_lnk_up = '0' then
      --if reset = '0' then
         rdndreqpipeline <= (others => '0');
      elsif rdndreqpipelineincr = '1' and rdndreqpipelinedecr = '1' then
         rdndreqpipeline <= rdndreqpipeline;
      elsif rdndreqpipelineincr = '1' then
         rdndreqpipeline <= rdndreqpipeline + 1;
      elsif rdndreqpipelinedecr = '1' then
         rdndreqpipeline <= rdndreqpipeline - 1;
      end if;
   end if;
end process;
end generate;

rd_req_128: if C_S_AXIS_DATA_WIDTH = 128 generate
rd_req_pipeline: process(aclk)
begin
   --pipeline buffer availability up/counter counter - CplD
   if rising_edge(aclk) then
      if reset = '0' or blk_lnk_up = '0' then
         rdreqpipeline <= (others => '0');
      elsif s_axis_cr_tvalid = '1' and s_axis_cr_tready_sig = '1' and rdreqpipelinedecr = '1' and s_axis_cr_tdata(30) = '0' and 
         s_axis_cr_tdata(28 downto 24) = "00000" and ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '1') or (C_PCIEBAR_NUM > 1 and
         ( s_axis_cr_tuser(2) = '1' or s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) and 
         s_axis_cr_tdata(35 downto 32) /= "0000" then
         rdreqpipeline <= rdreqpipeline;
      elsif s_axis_cr_tvalid = '1' and s_axis_cr_tready_sig = '1' and s_axis_cr_tdata(30) = '0' and 
         s_axis_cr_tdata(28 downto 24) = "00000" and ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '1') or (C_PCIEBAR_NUM > 1 and
         ( s_axis_cr_tuser(2) = '1' or s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) and 
         s_axis_cr_tdata(35 downto 32) /= "0000" then
         rdreqpipeline <= rdreqpipeline + 1;
      elsif rdreqpipelinedecr = '1' then
         rdreqpipeline <= rdreqpipeline - 1;
      end if;
   end if;
   --pipeline buffer availability up/counter counter - Cpl
   if rising_edge(aclk) then
      if reset = '0' or blk_lnk_up = '0' then
         rdndreqpipeline <= (others => '0');
      elsif s_axis_cr_tvalid = '1' and s_axis_cr_tready_sig = '1' and rdndreqpipelinedecr = '1' and s_axis_cr_tdata(30) = '0' and 
         s_axis_cr_tdata(28 downto 24) = "00000" and ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '0') or (C_PCIEBAR_NUM > 1 and 
         s_axis_cr_tuser(2) = '0' and s_axis_cr_tuser(3) = '0' and s_axis_cr_tuser(4) = '0' and s_axis_cr_tuser(6) = '0')) then
         rdndreqpipeline <= rdndreqpipeline;
      elsif s_axis_cr_tvalid = '1' and s_axis_cr_tready_sig = '1' and rdndreqpipelinedecr = '1' and s_axis_cr_tdata(30) = '0' and 
         s_axis_cr_tdata(28 downto 24) = "00000" and ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '1') or (C_PCIEBAR_NUM > 1 and 
         ( s_axis_cr_tuser(2) = '1' or s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) and 
         s_axis_cr_tdata(35 downto 32) = "0000" then
         rdndreqpipeline <= rdndreqpipeline;
      elsif s_axis_cr_tvalid = '1' and s_axis_cr_tready_sig = '1' and s_axis_cr_tdata(30) = '0' and 
         s_axis_cr_tdata(28 downto 24) = "00000" and ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '0') or (C_PCIEBAR_NUM > 1 and 
         s_axis_cr_tuser(2) = '0' and s_axis_cr_tuser(3) = '0' and s_axis_cr_tuser(4) = '0' and s_axis_cr_tuser(6) = '0')) then
         rdndreqpipeline <= rdndreqpipeline + 1;
      elsif s_axis_cr_tvalid = '1' and s_axis_cr_tready_sig = '1' and s_axis_cr_tdata(30) = '0' and 
         s_axis_cr_tdata(28 downto 24) = "00000" and ((C_PCIEBAR_NUM = 1 and s_axis_cr_tuser(2) = '1') or (C_PCIEBAR_NUM > 1 and 
         (s_axis_cr_tuser(2) = '1' or s_axis_cr_tuser(3) = '1' or s_axis_cr_tuser(4) = '1' or s_axis_cr_tuser(6) = '1'))) and
         s_axis_cr_tdata(35 downto 32) = "0000" then
         rdndreqpipeline <= rdndreqpipeline + 1;
      elsif rdndreqpipelinedecr = '1' then
         rdndreqpipeline <= rdndreqpipeline - 1;
      end if;
   end if;
end process;
end generate;

cpld_packet_split: process(aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         ctargetpipeline <= (others => '0');
         length_offset <= (others => '0');
         cpldsplitsm <= idle;
      else
      case cpldsplitsm is
      --count calculation for # of compl per read req
         when idle =>
            if ctargetpipeline /= rdtargetpipeline then
               cpldsplitsm <= cpldsplitcalc;
               case blk_dcontrol(7 downto 5) is 
                  when "000" =>
                     if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                        length_offset(11 downto 2) <= (tlplength(conv_integer(ctargetpipeline(1 downto 0))) + 
                           tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(6 downto 2)) - 1;
                     else
                        length_offset <= (others => '1');
                     end if;
                  
                  when "001" =>
                     if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                        length_offset(11 downto 2) <= (tlplength(conv_integer(ctargetpipeline(1 downto 0))) + 
                           tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(7 downto 2)) - 1;
                     else
                        length_offset <= (others => '1');
                     end if;
                  
                  -- coverage off
                  when "010" =>
                     if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                        length_offset(11 downto 2) <= (tlplength(conv_integer(ctargetpipeline(1 downto 0))) + 
                           tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(8 downto 2)) - 1;
                     else
                        length_offset <= (others => '1');
                     end if;
                  
                  when "011" =>
                     if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                        length_offset(11 downto 2) <= (tlplength(conv_integer(ctargetpipeline(1 downto 0))) + 
                           tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(9 downto 2)) - 1;
                     else
                        length_offset <= (others => '1');
                     end if;
                  
                  when "100" =>
                     if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                        length_offset(11 downto 2) <= (tlplength(conv_integer(ctargetpipeline(1 downto 0))) + 
                           tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(10 downto 2)) - 1;
                     else
                        length_offset <= (others => '1');
                     end if;
                  
                  when "101" =>
                     if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                        length_offset(11 downto 2) <= (tlplength(conv_integer(ctargetpipeline(1 downto 0))) + 
                           tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(11 downto 2)) - 1;
                     else
                        length_offset <= (others => '1');
                     end if;
                  
                  when others =>
                     cpldsplitsm <= idle;
                  -- coverage on
               end case;
            else
               cpldsplitsm <= idle;
            end if;
         
         when cpldsplitcalc =>
            cpldsplitsm <= cpldsplitparam;
            case blk_dcontrol(7 downto 5) is 
               when "000" =>
                  if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                     if conv_integer(tlplength(conv_integer(ctargetpipeline(1 downto 0)))) > 32 then
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= length_offset(11 downto 7);
                     else
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00000";
                     end if;
                  else
                     cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "11111";
                  end if;
               
               when "001" =>
                  if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                     if conv_integer(tlplength(conv_integer(ctargetpipeline(1 downto 0)))) > 64 then
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= '0' & length_offset(11 downto 8);
                     else
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00000";
                     end if;
                  else
                     cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "01111";
                  end if;
               
               -- coverage off
               when "010" =>
                  if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                     if conv_integer(tlplength(conv_integer(ctargetpipeline(1 downto 0)))) > 128 then
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00" & length_offset(11 downto 9);
                     else
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00000";
                     end if;
                  else
                     cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00111";
                  end if;
               
               when "011" =>
                  if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                     if conv_integer(tlplength(conv_integer(ctargetpipeline(1 downto 0)))) > 256 then
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "000" & length_offset(11 downto 10);
                     else
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00000";
                     end if;
                  else
                     cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00011";
                  end if;
               
               when "100" =>
                  if tlplength(conv_integer(ctargetpipeline(1 downto 0))) /= "0000000000" then
                     if conv_integer(tlplength(conv_integer(ctargetpipeline(1 downto 0)))) > 512 then
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "0000" & length_offset(11 downto 11);
                     else
                        cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00000";
                     end if;
                  else
                     cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00001";
                  end if;
               
               when "101" =>
                  cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0))) <= "00000";
               
               when others =>
                  cpldsplitsm <= idle;
               -- coverage on
            end case;
         
         when cpldsplitparam =>
         --completion splits header info (len, bytecount)
            case blk_dcontrol(7 downto 5) is 
               when "000" =>
                  if conv_integer(cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0)))) = 0 then
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                        tlplength(conv_integer(ctargetpipeline(1 downto 0)));
                  else
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & x"20" - 
                        tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(6 downto 2);
                  end if;
                  ctlplength(1, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & x"20";
                  ctlplength(2, conv_integer(ctargetpipeline(1 downto 0))) <= "00000" & length_offset(6 downto 2) + 1;
                  ctlpbytecount(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlpbytecount(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlpbytecount(1, conv_integer(ctargetpipeline(1 downto 0))) <= x"080" - 
                     tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(6 downto 0);
               
               when "001" =>
                  if conv_integer(cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0)))) = 0 then
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                        tlplength(conv_integer(ctargetpipeline(1 downto 0)));
                  else
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & x"40" - 
                        tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(7 downto 2);
                  end if;
                  ctlplength(1, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & x"40";
                  ctlplength(2, conv_integer(ctargetpipeline(1 downto 0))) <= "0000" & length_offset(7 downto 2) + 1;
                  ctlpbytecount(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlpbytecount(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlpbytecount(1, conv_integer(ctargetpipeline(1 downto 0))) <= x"100" - 
                     tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(7 downto 0);
               
               -- coverage off
               when "010" =>
                  if conv_integer(cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0)))) = 0 then
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                        tlplength(conv_integer(ctargetpipeline(1 downto 0)));
                  else
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & x"80" - 
                        tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(8 downto 2);
                  end if;
                  ctlplength(1, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & x"80";
                  ctlplength(2, conv_integer(ctargetpipeline(1 downto 0))) <= "000" & length_offset(8 downto 2) + 1;
                  ctlpbytecount(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlpbytecount(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlpbytecount(1, conv_integer(ctargetpipeline(1 downto 0))) <= x"200" - 
                     tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(8 downto 0);
               
               when "011" =>
                  if conv_integer(cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0)))) = 0 then
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                        tlplength(conv_integer(ctargetpipeline(1 downto 0)));
                  else
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= "01" & x"00" - 
                        tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(9 downto 2);
                  end if;
                  ctlplength(1, conv_integer(ctargetpipeline(1 downto 0))) <= "01" & x"00";
                  ctlplength(2, conv_integer(ctargetpipeline(1 downto 0))) <= "00" & length_offset(9 downto 2) + 1;
                  ctlpbytecount(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlpbytecount(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlpbytecount(1, conv_integer(ctargetpipeline(1 downto 0))) <= x"400" - 
                     tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(9 downto 0);
               
               when "100" =>
                  if conv_integer(cpldsplitcount(conv_integer(ctargetpipeline(1 downto 0)))) = 0 then
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                        tlplength(conv_integer(ctargetpipeline(1 downto 0)));
                  else
                     ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= "10" & x"00" - 
                        tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(10 downto 2);
                  end if;
                  ctlplength(1, conv_integer(ctargetpipeline(1 downto 0))) <= (others => '0');
                  ctlplength(2, conv_integer(ctargetpipeline(1 downto 0))) <= '0' & length_offset(10 downto 2) + 1;
                  ctlpbytecount(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlpbytecount(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlpbytecount(1, conv_integer(ctargetpipeline(1 downto 0))) <= x"800" - 
                     tlpaddrl(conv_integer(ctargetpipeline(1 downto 0)))(10 downto 0);
               
               when "101" =>
                  ctlplength(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlplength(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlplength(1, conv_integer(ctargetpipeline(1 downto 0))) <= (others => '0');
                  ctlplength(2, conv_integer(ctargetpipeline(1 downto 0))) <= (others => '0');
                  ctlpbytecount(0, conv_integer(ctargetpipeline(1 downto 0))) <= 
                     tlpbytecount(conv_integer(ctargetpipeline(1 downto 0)));
                  ctlpbytecount(1, conv_integer(ctargetpipeline(1 downto 0))) <= (others => '0');
               
               when others =>
                  cpldsplitsm <= idle;
               -- coverage on
            end case;
            ctargetpipeline <= ctargetpipeline + 1;
            cpldsplitsm <= idle;
            
         -- coverage off
         when others =>
            cpldsplitsm <= idle;
         -- coverage on
      end case;
      if blk_lnk_up_latch = '0' and cpltargetpipeline /= ctargetpipeline then
         ctargetpipeline <= addrstreampipeline;
      end if;
      end if;
   end if;
end process;

m_axis_cc_tvalid <= m_axis_cc_tvalid_nd when cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline else
                    m_axis_cc_tvalid_d;
dw32: if C_S_AXIS_DATA_WIDTH = 32 generate
m_axis_cc_tdata_d <= m_axis_cc_tdata_h when data_phase = '0' else
                     little_to_big_endian32(dout);
end generate dw32;

dw64: if C_S_AXIS_DATA_WIDTH = 64 generate
m_axis_cc_tdata_d <= m_axis_cc_tdata_h when data_phase = '0' else
                     little_to_big_endian32(dout(63 downto 32)) & little_to_big_endian32(dout(31 downto 0)) 
                        when (cplpacket1 = '1' and rdtlpaddrltemp(2) = '1') else
                     little_to_big_endian32(dout(31 downto 0)) & little_to_big_endian32(m_axis_cc_tdatatemp64);
end generate dw64;

dw128: if C_S_AXIS_DATA_WIDTH = 128 generate
m_axis_cc_tdata_d <= m_axis_cc_tdata_h when data_phase = '0' else
                     little_to_big_endian32(dout(127 downto 96)) & little_to_big_endian32(dout(95 downto 64)) & 
                        little_to_big_endian32(dout(63 downto 32)) & little_to_big_endian32(dout(31 downto 0)) 
                           when cplpacket1 = '1' and rdtlpaddrltemp(3 downto 2) = "11" else
                     little_to_big_endian32(dout(95 downto 64)) & little_to_big_endian32(dout(63 downto 32)) & 
                        little_to_big_endian32(dout(31 downto 0)) & little_to_big_endian32(m_axis_cc_tdatatemp128(95 downto 64)) 
                           when cplpacket1 = '1' and rdtlpaddrltemp(3) = '1' else
                     little_to_big_endian32(dout(63 downto 32)) & little_to_big_endian32(dout(31 downto 0)) & 
                        little_to_big_endian32(m_axis_cc_tdatatemp128(95 downto 64)) & 
                           little_to_big_endian32(m_axis_cc_tdatatemp128(63 downto 32)) 
                              when cplpacket1 = '1' and rdtlpaddrltemp(2) = '1' else
                     little_to_big_endian32(dout(31 downto 0)) & little_to_big_endian32(m_axis_cc_tdatatemp128(95 downto 64)) & 
                        little_to_big_endian32(m_axis_cc_tdatatemp128(63 downto 32)) & 
                           little_to_big_endian32(m_axis_cc_tdatatemp128(31 downto 0));
end generate dw128;

-- modified rd_en expression, CR #671086 (AXI PCIE 37x BURST ISSUE)

rd_en64_32: if C_S_AXIS_DATA_WIDTH /= 128 generate
rd_en            <= (m_axis_cc_tready or corruptdataflush or lnkdowndataflush) and (m_axis_cc_tvalid_d or rd_en_sig) and 
                       not(empty) and (data_phase or rd_en_sig) and not(dis_rden);
end generate rd_en64_32;

rd_en128: if C_S_AXIS_DATA_WIDTH = 128 generate
rd_en            <= (rd_en_sig or m_axis_cc_tready or corruptdataflush or lnkdowndataflush) and (m_axis_cc_tvalid_d or rd_en_sig) and 
                       		not(empty) and (data_phase or rd_en_sig) and not(dis_rden) when (cpltlpsmsig = memcpltxonedw or (cpltlpsmsig = memcpltxdata and ctlplengthtemp = "0000000001")) else
                    (m_axis_cc_tready or corruptdataflush or lnkdowndataflush) and (m_axis_cc_tvalid_d or rd_en_sig) and 
                       		not(empty) and (data_phase or rd_en_sig) and not(dis_rden);
end generate rd_en128;


m_axis_cc_tdata <= m_axis_cc_tdata_nd when cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline else
                   m_axis_cc_tdata_d;
m_axis_cc_tstrb <= m_axis_cc_tstrb_nd when cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline else
                   m_axis_cc_tstrb_d;
m_axis_cc_tlast <= m_axis_cc_tlast_nd when cplndtargetpipeline /= rdndtargetpipeline and cpltlpsmsig = memcplpipeline else
                   m_axis_cc_tlast_d;

rdtargetpipeline_out <= rdtargetpipeline;

s_axis_cr_tready <= s_axis_cr_tready_sig;

m_axis_cc_tuser <= (others => '0');

wrpending <= wrpendingsig;

end behavioral;




-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_s_masterbridge_wr.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge write function
-- on the AXI Stream.
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_s_masterbridge_wr.vhd
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

--library AMDCoreLib;
--use AMDCoreLib.all;
--library UNISIM;
--use UNISIM.VComponents.all;

entity axi_s_masterbridge_wr is
   generic(
      --Family Generics
      C_FAMILY            : string;
      C_S_AXIS_DATA_WIDTH : integer;
      C_S_AXIS_USER_WIDTH : integer;
      C_PCIEBAR_NUM       : integer
      );
   port(
      --AXI Global
      aclk             : in  std_logic; --meaningful port name
      reset            : in  std_logic; --meaningful port name
      --AXIS Write Target Channel
      s_axis_cw_tdata  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      s_axis_cw_tstrb  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name (not used)
      s_axis_cw_tlast  : in  std_logic; --meaningful port name
      s_axis_cw_tvalid : in  std_logic; --meaningful port name
      s_axis_cw_tready : out std_logic; --meaningful port name
      s_axis_cw_tuser  : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --Master Bridge Interrupt Strobes
      master_int       : out std_logic; --meaningful port name
      --AXI Streaming Block Interface
      blk_lnk_up       : in  std_logic; --meaningful port name
      --Internal Interface
      tlplength          : out std_logic_vector(9 downto 0); --meaningful port name
      firstdwbe          : out std_logic_vector(3 downto 0); --meaningful port name
      lastdwbe           : out std_logic_vector(3 downto 0); --meaningful port name
      tlpaddrl           : out std_logic_vector(31 downto 0); --meaningful port name
      tlpaddrh           : out std_logic_vector(31 downto 0); --meaningful port name
      datain             : out std_logic_vector(C_S_AXIS_DATA_WIDTH downto 0); --meaningful port name
      wrreqset           : out std_logic; --meaningful port name
      datacompcheck      : in  std_logic; --meaningful port name (used for testing)
      tlppipeline        : in  std_logic_vector(2 downto 0); --meaningful port name
      dataen             : out std_logic; --meaningful port name
      almost_full        : in  std_logic; --meaningful port name
      wrreqpend          : out std_logic_vector(2 downto 0); --meaningful port name
      treadydataenadjust : out std_logic --meaningful port name
      );
end axi_s_masterbridge_wr;

architecture behavioral of axi_s_masterbridge_wr is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

type wr_master_ingress_states is (idle,
                                  memwrreq,
                                  onedwlength,
                                  zerolenwr,
                                  poisoneddataclkout,
                                  blklinkdown,
                                  throttle,
                                  latchbe,
                                  latchaddrh,
                                  latchaddrl,
                                  datatransfer);

signal wrreqsmsig                            : wr_master_ingress_states;
signal wrreqsetsig                           : std_logic;
signal tlpepsig                              : std_logic;
signal tlpfmtsig                             : std_logic_vector(1 downto 0);
signal tlptypesig                            : std_logic_vector(4 downto 0);
signal tlplengthsig                          : std_logic_vector(9 downto 0);
signal firstdwbesig, lastdwbesig             : std_logic_vector(3 downto 0);
signal delaylast,  s_axis_cw_tlasttemp       : std_logic;
signal tempdatareg                           : std_logic_vector(31 downto 0);
signal s_axis_cw_tdatatemp                   : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
signal dataoffset, addroffset                : std_logic;
signal addroffset1, addroffset2, addroffset3 : std_logic;
signal padzeroes                             : std_logic;
signal blk_lnk_upsig                         : std_logic;
signal s_axis_cw_treadysig                   : std_logic;
signal wrreqpendsig                          : std_logic_vector(2 downto 0);

function little_to_big_endian32(datain : std_logic_vector(31 downto 0))
      return std_logic_vector is
   variable dataout : std_logic_vector(31 downto 0);
begin
   dataout := datain(7 downto 0) & datain(15 downto 8) & datain(23 downto 16) & datain(31 downto 24);
   return(dataout);
end function;

begin

data_width_32: if C_S_AXIS_DATA_WIDTH = 32 generate
wr_master_ingress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cw_treadysig    <= '0';
         tlplengthsig        <= (others => '0');
         firstdwbesig        <= (others => '0');
         lastdwbesig         <= (others => '0');
         tlpaddrl            <= (others => '0');
         tlpaddrh            <= (others => '0');
         tlpfmtsig           <= (others => '0');
         tlptypesig          <= (others => '0');
         s_axis_cw_tdatatemp <= (others => '0');
         dataen              <= '0';
         wrreqsmsig          <= idle;
         datain              <= (others => '0');
         wrreqsetsig         <= '0';
         master_int          <= '0';
         delaylast           <= '0';
         dataoffset          <= '0';
         addroffset          <= '0';
         addroffset1         <= '0';
         addroffset2         <= '0';
         addroffset3         <= '0';
         padzeroes           <= '0';
         s_axis_cw_tlasttemp <= '0';
         tempdatareg         <= (others => '0');
         blk_lnk_upsig       <= '0';
         wrreqpendsig        <= "000";
      else
         case wrreqsmsig is
            when idle =>
               if tlppipeline /= "100" then
                  s_axis_cw_treadysig <= '1';
                  wrreqsmsig       <= memwrreq;
               end if;
               tlplengthsig     <= (others => '0');
               firstdwbesig     <= (others => '0');
               lastdwbesig      <= (others => '0');
               tlpaddrl         <= (others => '0');
               tlpaddrh         <= (others => '0');
               tlpfmtsig        <= (others => '0');
               tlptypesig       <= (others => '0');
               dataen           <= '0';
               datain           <= (others => '0');
               wrreqsetsig      <= '0';
               master_int       <= '0';
               blk_lnk_upsig    <= '0';

           
            when memwrreq=>
               -- Nam -- extremely hard to hit case for FALSE branch
               -- NAM / JRH fixed typo. Was b 2.
               -- coverage off -item b 1 -allfalse
               if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     tlpepsig <= s_axis_cw_tdata(14);
                  -- Nam - double check
                  -- coverage off -item b 1 -allfalse                            
                     if s_axis_cw_tdata(30) = '1' then
                        -- Nam - -- tool issue, work work when the if statement is more than 1 line
                        -- coverage off -item bc 1 -allfalse -condrow 1 2 6
                        if s_axis_cw_tdata(28 downto 24) = "00000" and (s_axis_cw_tuser(2) = '1' or 
                           s_axis_cw_tuser(3) = '1' or s_axis_cw_tuser(4) = '1' or s_axis_cw_tuser(6) = '1') then
                           if s_axis_cw_tdata(14) = '0' then
                              tlpfmtsig    <= s_axis_cw_tdata(30 downto 29);
                              tlptypesig   <= s_axis_cw_tdata(28 downto 24);
                              tlplengthsig <= s_axis_cw_tdata(9 downto 0);
                              wrreqsmsig   <= latchbe;
                           else
                              wrreqsmsig    <= poisoneddataclkout;
                              master_int <= '1';
                           end if;
                        end if;
                     end if;
                  end if;
               end if;

            when poisoneddataclkout =>
               master_int <= '0';
               if blk_lnk_up = '1' then
                  -- Nam - enhance bridge wont throttle
                  -- coverage off -item b 1 -allfalse                      
                  if s_axis_cw_tvalid = '1' then
                     if s_axis_cw_tlast = '1' then
                        wrreqsmsig       <= memwrreq;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - poison data while linkdown
               -- coverage off
               else
                  if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                     wrreqsmsig       <= memwrreq;
                  else
                     wrreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            
            when blklinkdown =>
               -- Nam - enhance bridge wont throttle
               -- coverage off -item b 1 -allfalse                
               if s_axis_cw_tvalid = '1' then
                  -- Nam - enhance bridge wont throttle
                  -- coverage off -item b 1 -allfalse                      
                  if s_axis_cw_tlast = '1' then
                     wrreqsmsig       <= idle;
                  end if;
               else
                  wrreqsmsig     <= idle;
               end if;
            
            when latchbe =>
               if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     if s_axis_cw_tdata(3 downto 0) /= "0000" then
                        lastdwbesig  <= s_axis_cw_tdata(7 downto 4);
                        firstdwbesig <= s_axis_cw_tdata(3 downto 0);
                        if tlpfmtsig(0) = '0' then
                           wrreqsmsig  <= latchaddrl;
                        else
                           wrreqsmsig <= latchaddrh;
                        end if;
                     else
                        wrreqsmsig       <= zerolenwr;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - we cover this with 2 hits during the weekend run
               -- coverage off                  
               else
                  wrreqsmsig       <= blklinkdown;
               end if;
               -- coverage on

            when zerolenwr =>
               if blk_lnk_up = '1' then
                   -- Nam - enhance bridge wont throttle
                   -- coverage off -item b 1 -allfalse                      
                   if s_axis_cw_tvalid = '1' then
                     if s_axis_cw_tlast = '1' then
                        s_axis_cw_treadysig <= '0';
                        wrreqsmsig       <= idle;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - zero length write while linkdown
               -- coverage off                  
               else
                  if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                     s_axis_cw_treadysig <= '0';
                     wrreqsmsig       <= idle;
                  else
                     wrreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            
            when latchaddrh =>
               if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     tlpaddrh    <= s_axis_cw_tdata;
                     wrreqsmsig  <= latchaddrl;
                  end if;
               -- Nam -- extremely hard to hit case - we cover this with 1 hits during the weekend run
               -- coverage off                   
               else
                  wrreqsmsig       <= blklinkdown;
               end if;
               -- coverage on
               
            when latchaddrl =>
               if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     if tlppipeline /= "100" then
                        wrreqsetsig <= '1';
                        wrreqpendsig <= wrreqpendsig + 1;
                        tlpaddrl <= s_axis_cw_tdata;
                        dataen <= '1';
                        wrreqsmsig <= datatransfer;
                     else
                        wrreqsmsig <= throttle;
                        s_axis_cw_treadysig <= '0';
                        tlpaddrl <= s_axis_cw_tdata;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - we cover this with 2 hits during the weekend run
               -- coverage off                   
               else
                  wrreqsmsig       <= blklinkdown;
               end if;
               -- coverage on
            when throttle =>
               if blk_lnk_up = '1' then
                  if tlppipeline /= "100" then
                     wrreqsetsig <= '1';
                     wrreqpendsig <= wrreqpendsig + 1;
                     dataen      <= '1';
                     wrreqsmsig   <= datatransfer;
                     s_axis_cw_treadysig <= '1';
                  end if;
               else
                  wrreqsmsig    <= blklinkdown;
                  s_axis_cw_treadysig <= '1';
               end if;

            when datatransfer =>
               wrreqsetsig <= '0';
               -- Nam - enhance core does not throttle
               -- coverage off -item b 1 -allfalse
               if s_axis_cw_tvalid = '1' then
                  s_axis_cw_treadysig <= not(almost_full);
                  if almost_full = '0' then
                     if s_axis_cw_treadysig = '1' then
                        dataen <= '1';
                        datain <= s_axis_cw_tlast & little_to_big_endian32(s_axis_cw_tdata);
                        if s_axis_cw_tlast = '1' then
                           wrreqsmsig <= idle;
                           dataen     <= '0';
                           s_axis_cw_treadysig <= '0';
                        end if;                                         
                     end if;
                  end if;
               end if;
               if blk_lnk_up = '0' then
                  blk_lnk_upsig <= '1';
               end if;


            -- coverage off
            when others => wrreqsmsig <= idle;
            -- coverage on
         end case;
      end if;
   end if;
end process;
end generate;

data_width_64: if C_S_AXIS_DATA_WIDTH = 64 generate
wr_master_ingress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cw_treadysig    <= '0';
         tlplengthsig        <= (others => '0');
         firstdwbesig        <= (others => '0');
         lastdwbesig         <= (others => '0');
         tlpaddrl            <= (others => '0');
         tlpaddrh            <= (others => '0');
         tlpfmtsig           <= (others => '0');
         tlptypesig          <= (others => '0');
         s_axis_cw_tdatatemp <= (others => '0');
         dataen              <= '0';
         wrreqsmsig          <= idle;
         datain              <= (others => '0');
         wrreqsetsig         <= '0';
         master_int          <= '0';
         delaylast           <= '0';
         dataoffset          <= '0';
         addroffset          <= '0';
         addroffset1         <= '0';
         addroffset2         <= '0';
         addroffset3         <= '0';
         padzeroes           <= '0';
         s_axis_cw_tlasttemp <= '0';
         tempdatareg         <= (others => '0');
         blk_lnk_upsig       <= '0';
         wrreqpendsig        <= "000";
      else
         case wrreqsmsig is
            when idle =>
               if tlppipeline /= "100" then
                  s_axis_cw_treadysig <= '1';
                  wrreqsmsig       <= memwrreq;
               end if;
               delaylast           <= '0';
               tlplengthsig        <= (others => '0');
               firstdwbesig        <= (others => '0');
               lastdwbesig         <= (others => '0');
               tlpaddrl            <= (others => '0');
               tlpaddrh            <= (others => '0');
               tlpfmtsig           <= (others => '0');
               tlptypesig          <= (others => '0');
               dataen              <= '0';
               datain              <= (others => '0');
               wrreqsetsig         <= '0';
               master_int          <= '0';
               blk_lnk_upsig       <= '0';
               dataoffset          <= '0';
               addroffset          <= '0';
               padzeroes           <= '0';
               s_axis_cw_tlasttemp <= '0';
               tempdatareg         <= (others => '0');

            
            when memwrreq =>
               wrreqsetsig <= '0';
               addroffset  <= '0';
               -- Nam -- extremely hard to hit case for FALSE branch
               -- NAM / JRH fixed typo. Was b 2.
               -- coverage off -item b 1 -allfalse
               if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     tlpepsig <= s_axis_cw_tdata(14);
                     -- Nam - double check
                     -- coverage off -item b 1 -allfalse
                     if s_axis_cw_tdata(30) = '1' then
                        -- Nam - -- tool issue, work work when the if statement is more than 1 line
                        -- coverage off -item bc 1 -allfalse -condrow 1 2 6
                        if s_axis_cw_tdata(28 downto 24) = "00000" and ((s_axis_cw_tuser(2) = '1' and C_PCIEBAR_NUM = 1)
                          or (C_PCIEBAR_NUM > 1 and (s_axis_cw_tuser(2) = '1' or s_axis_cw_tuser(3) = '1' or 
                          s_axis_cw_tuser(4) = '1' or s_axis_cw_tuser(6) = '1'))) then
                           if s_axis_cw_tdata(14) = '0' then
                              tlpfmtsig     <= s_axis_cw_tdata(30 downto 29);
                              tlptypesig    <= s_axis_cw_tdata(28 downto 24);
                              tlplengthsig  <= s_axis_cw_tdata(9 downto 0);
                              lastdwbesig   <= s_axis_cw_tdata(39 downto 36);
                              firstdwbesig  <= s_axis_cw_tdata(35 downto 32);
                              if s_axis_cw_tdata(35 downto 32) /= "0000" then
                                 if wrreqsetsig = '0' and tlppipeline /= "100" then
                                    if s_axis_cw_tdata(29) = '0' then
                                       wrreqsmsig <= latchaddrl;
                                       if s_axis_cw_tdata(9 downto 0) = 1 then
                                          dataen  <= '1';
                                       end if;
                                    else
                                       wrreqsmsig <= latchaddrh;
                                    end if;
                                 else
                                    wrreqsmsig    <= throttle;
                                    s_axis_cw_treadysig <= '0';
                                 end if;
                              else
                                 wrreqsmsig       <= zerolenwr;
                              end if;
                           else
                              wrreqsmsig    <= poisoneddataclkout;
                              master_int <= '1';
                           end if;
                        end if;
                     end if;
                  end if;
                  blk_lnk_upsig  <= '0';
               end if;
            
            when poisoneddataclkout =>
               s_axis_cw_treadysig <= s_axis_cw_treadysig;
	       master_int <= '0';
               if blk_lnk_up = '1' then
                  -- Nam - enhance bridge wont throttle
                  -- coverage off -item b 1 -allfalse
                  if s_axis_cw_tvalid = '1' then
                     if s_axis_cw_tlast = '1' then
                        wrreqsmsig       <= memwrreq;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - poison data while linkdown
               -- coverage off                  
               else
                  if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                     wrreqsmsig       <= memwrreq;
                  else
                     wrreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            
            when blklinkdown =>
	       s_axis_cw_treadysig <= s_axis_cw_treadysig;
               -- Nam - enhance bridge wont throttle
               -- coverage off -item b 1 -allfalse            
               if s_axis_cw_tvalid = '1' then
                  if s_axis_cw_tlast = '1' then
                     wrreqsmsig     <= idle;
                  end if;
               else
                  wrreqsmsig     <= idle;
               end if;
            
            when zerolenwr =>
               if blk_lnk_up = '1' then
                  -- Nam - enhance core does not throttle
                  -- coverage off -item b 1 -allfalse
                  if s_axis_cw_tvalid = '1' then
                     if s_axis_cw_tlast = '1' then
                        s_axis_cw_treadysig <= '0';
                        wrreqsmsig       <= idle;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - zero length write while link_down
               -- coverage off
               else
                   if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                      s_axis_cw_treadysig <= '0';
                      wrreqsmsig       <= idle;
                   else
                      wrreqsmsig       <= blklinkdown;
                   end if;
               end if;
               -- coverage on

            when throttle =>
               if blk_lnk_up = '1' then
                  if tlppipeline /= "100" then
                     s_axis_cw_treadysig <= '1';
                     if tlpfmtsig(0) = '0' then
                        wrreqsmsig    <= latchaddrl;
                        if s_axis_cw_tlast = '1' then
                           dataen     <= '1';
                        end if;
                     else
                        wrreqsmsig   <= latchaddrh;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case. We covered this with the weekend run - 10 hits
               -- coverage off
               else
                  wrreqsmsig    <= blklinkdown;
                  s_axis_cw_treadysig <= '1';
               end if;
               -- coverage on
               
            when latchaddrh =>
               s_axis_cw_treadysig <= s_axis_cw_treadysig;
	       if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     wrreqsetsig <= '1';
                     wrreqpendsig <= wrreqpendsig + 1;
                     tlpaddrh    <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 0);
                     tlpaddrl    <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto C_S_AXIS_DATA_WIDTH/2);
                     if s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) = '1' then
                        addroffset   <= '1';
                        padzeroes    <= '1';
                        if tlplengthsig(0) = '0' then
                           delaylast <= '1';
                        end if;
                     end if;
                     dataen     <= '1';
                     wrreqsmsig <= datatransfer;
                  end if;
               -- Nam -- extremely hard to hit case. We covered this with the weekend run - 2 hits
               -- coverage off                  
               else
                  wrreqsmsig    <= blklinkdown;
               end if;
               -- coverage on

            when latchaddrl =>
               s_axis_cw_treadysig <= s_axis_cw_treadysig;
	       if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     wrreqsetsig <= '1';
                     wrreqpendsig <= wrreqpendsig + 1;
                     tlpaddrl    <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 0);
                     if s_axis_cw_tdata(2) = '1' then
                        addroffset   <= '1';
                        if s_axis_cw_tlast = '0' then
                           padzeroes <= '1';
                        end if;
                     end if;
                     tempdatareg <= little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto C_S_AXIS_DATA_WIDTH/2));
                     if s_axis_cw_tlast = '1' then
                        if s_axis_cw_tdata(2) = '1' then
                           datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto C_S_AXIS_DATA_WIDTH/2)) & 
                                x"0000_0000";
                        else
                           datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= x"0000_0000" & 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto C_S_AXIS_DATA_WIDTH/2));
                        end if;
                        datain(C_S_AXIS_DATA_WIDTH)  <= '1';
                        wrreqsmsig <= memwrreq;
                        dataen     <= '0';
                     else
                        dataoffset   <= '1';
                        dataen       <= '1';
                        wrreqsmsig   <= datatransfer;
                        if tlplengthsig(0) = '1' or s_axis_cw_tdata(2) = '1' then
                           delaylast <= '1';
                        end if;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case.  
               -- coverage off                  
               else
                  if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                     wrreqsmsig       <= idle;
                  else
                     wrreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on

            when datatransfer =>
               wrreqsetsig <= '0';
               -- Nam - enhance bridge wont throttle -  -- tool issue, work work when the if statement is more than 1 line
               -- coverage off -item bc 1 -allfalse -condrow 3
               if s_axis_cw_tvalid = '1' or s_axis_cw_tlasttemp = '1' then
                  s_axis_cw_treadysig <= not(almost_full);
                  if almost_full = '0' then
                  if s_axis_cw_treadysig = '1' or s_axis_cw_tlasttemp = '1' then
                  if dataoffset  = '1' then
                     if addroffset = '0' then
                        datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                          little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 0)) & 
                           tempdatareg;
                        tempdatareg <= little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto C_S_AXIS_DATA_WIDTH/2));
                     else
                        if padzeroes = '0' then
                           datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= s_axis_cw_tdatatemp;
                        else
                           datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= tempdatareg & x"00000000";
                           padzeroes <= '0';
                        end if;
                        s_axis_cw_tdatatemp <= little_to_big_endian32(s_axis_cw_tdata(63 downto 32)) & 
                          little_to_big_endian32(s_axis_cw_tdata(31 downto 0));
                     end if;
                  else
                     if addroffset = '0' then
                        datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= little_to_big_endian32(s_axis_cw_tdata(63 downto 32)) & 
                          little_to_big_endian32(s_axis_cw_tdata(31 downto 0));
                     else
                        if padzeroes = '0' then
                           datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                             little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 0)) 
                              & s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2-1 downto 0);
                        else
                           datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                             little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 0)) 
                              & x"00000000";
                           padzeroes <= '0';
                        end if;
                        s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2-1 downto 0) <= 
                           little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto C_S_AXIS_DATA_WIDTH/2));
                     end if;
                  end if;
                  if delaylast = '0' then
                     datain(C_S_AXIS_DATA_WIDTH) <= s_axis_cw_tlast;
                     if s_axis_cw_tlast = '1' then
                        s_axis_cw_treadysig <= '0';
                        wrreqsmsig <= idle;
                        dataen     <= '0';
                        dataoffset <= '0';
                        addroffset <= '0';
                     end if;
                  else
                     s_axis_cw_tlasttemp <= s_axis_cw_tlast;
                     datain(C_S_AXIS_DATA_WIDTH) <= s_axis_cw_tlasttemp;
                     if s_axis_cw_tlast = '1' then
                        s_axis_cw_treadysig <= '0';
                     end if;
                     if s_axis_cw_tlasttemp = '1' then
                        s_axis_cw_treadysig <= '0';
                        wrreqsmsig <= idle;
                        dataen     <= '0';
                        dataoffset <= '0';
                        delaylast  <= '0';
                        addroffset <= '0';
                        s_axis_cw_tlasttemp <= '0';
                     end if;
                  end if;
                  end if;
                  end if;
               end if;
               if blk_lnk_up = '0' then
                  blk_lnk_upsig <= '1';
               end if;

            -- coverage off
            when others =>
               s_axis_cw_treadysig <= s_axis_cw_treadysig;
	       wrreqsmsig <= idle;
            -- coverage on
         end case;
      end if;
   end if;
end process;
end generate;

data_width_128: if C_S_AXIS_DATA_WIDTH = 128 generate
wr_master_ingress: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cw_treadysig    <= '0';
         tlplengthsig        <= (others => '0');
         firstdwbesig        <= (others => '0');
         lastdwbesig         <= (others => '0');
         tlpaddrl            <= (others => '0');
         tlpaddrh            <= (others => '0');
         tlpfmtsig           <= (others => '0');
         tlptypesig          <= (others => '0');
         s_axis_cw_tdatatemp <= (others => '0');
         dataen              <= '0';
         wrreqsmsig          <= idle;
         datain              <= (others => '0');
         wrreqsetsig         <= '0';
         master_int          <= '0';
         delaylast           <= '0';
         dataoffset          <= '0';
         addroffset          <= '0';
         addroffset1         <= '0';
         addroffset2         <= '0';
         addroffset3         <= '0';
         padzeroes           <= '0';
         s_axis_cw_tlasttemp <= '0';
         tempdatareg         <= (others => '0');
         blk_lnk_upsig       <= '0';
         wrreqpendsig        <= "000";
      else
         case wrreqsmsig is
            when idle =>
               s_axis_cw_treadysig <= '1';
               delaylast <= '0';
               tlplengthsig     <= (others => '0');
               firstdwbesig     <= (others => '0');
               lastdwbesig      <= (others => '0');
               tlpaddrl         <= (others => '0');
               tlpaddrh         <= (others => '0');
               tlpfmtsig        <= (others => '0');
               tlptypesig       <= (others => '0');
               dataen           <= '0';
               wrreqsmsig       <= memwrreq;
               datain           <= (others => '0');
               wrreqsetsig      <= '0';
               master_int       <= '0';
               blk_lnk_upsig    <= '0';
               dataoffset       <= '0';
               addroffset1      <= '0';
               addroffset2      <= '0';
               addroffset3      <= '0';
               padzeroes        <= '0';
               s_axis_cw_tlasttemp <= '0';
               tempdatareg      <= (others => '0');

            
            when memwrreq =>
               -- Nam -- extremely hard to hit case for FALSE branch
               -- NAM / JRH fixed typo. Was b 2.
               -- coverage off -item b 1 -allfalse
               if blk_lnk_up = '1' then
                  if s_axis_cw_tvalid = '1' and almost_full = '0' then
                     tlpepsig <= s_axis_cw_tdata(14);
                     -- Nam - double check
                     -- coverage off -item b 1 -allfalse
                     if s_axis_cw_tdata(30) = '1' then
                        -- Nam - -- tool issue, work work when the if statement is more than 1 line
                        -- coverage off -item bc 1 -allfalse -condrow 1 2 6
                        if s_axis_cw_tdata(28 downto 24) = "00000" and ((s_axis_cw_tuser(2) = '1' and C_PCIEBAR_NUM = 1)
                          or (C_PCIEBAR_NUM > 1 and (s_axis_cw_tuser(2) = '1' or s_axis_cw_tuser(3) = '1' or 
                          s_axis_cw_tuser(4) = '1' or s_axis_cw_tuser(6) = '1'))) then
                           if s_axis_cw_tdata(14) = '0' then
                              tlpfmtsig     <= s_axis_cw_tdata(30 downto 29);
                              tlptypesig    <= s_axis_cw_tdata(28 downto 24);
                              tlplengthsig  <= s_axis_cw_tdata(9 downto 0);
                              lastdwbesig   <= s_axis_cw_tdata(39 downto 36);
                              firstdwbesig  <= s_axis_cw_tdata(35 downto 32);
                              if s_axis_cw_tdata(35 downto 32) /= "0000" then
                                 s_axis_cw_tlasttemp <= s_axis_cw_tlast;
                                 if s_axis_cw_tdata(29) = '0' then
                                    tlpaddrl    <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto
                                       C_S_AXIS_DATA_WIDTH/2);
                                    tempdatareg <= little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                       C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4));
                                 else
                                    tlpaddrh    <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto
                                       C_S_AXIS_DATA_WIDTH/2);
                                    tlpaddrl    <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                       C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4);
                                 end if;
                                 if s_axis_cw_tdata(29) = '1' then
                                    if s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2) = '1' or 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3) = '1' then
                                       addroffset1  <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2) 
                                          and not(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3));
                                       addroffset2  <= 
                                          not(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2)) and 
                                             s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3);
                                       addroffset3  <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2) 
                                          and s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3);
                                       padzeroes    <= '1';
                                    end if;
                                    if s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2) = '1' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3) = '0' and 
                                          s_axis_cw_tdata(1 downto 0) = "00" then
                                       delaylast         <= '1';
                                    elsif s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2) = '0' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3) = '1' and 
                                          (s_axis_cw_tdata(1 downto 0) = "00" or 
                                             s_axis_cw_tdata(1 downto 0) = "11") then
                                       delaylast         <= '1';
                                    elsif s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+2) = '1' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4+3) = '1' and 
                                          s_axis_cw_tdata(1 downto 0) /= "01" then
                                       delaylast         <= '1';
                                    end if;
                                 else
                                    if s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) = '1' or 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3) = '1' then
                                       addroffset1  <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) and 
                                          not(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3));
                                       addroffset2  <= not(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2)) and 
                                          s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3);
                                       addroffset3  <= s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) and 
                                          s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3);
                                       padzeroes    <= '1';
                                    end if;
                                    if s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) = '0' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3) = '0' and 
                                          s_axis_cw_tdata(1 downto 0) = "01" then
                                       delaylast         <= '1';
                                    elsif s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) = '1' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3) = '0' and 
                                          (s_axis_cw_tdata(1 downto 0) = "00" or 
                                             s_axis_cw_tdata(1 downto 0) = "01") then
                                       delaylast         <= '1';
                                    elsif s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) = '0' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3) = '1' and 
                                          s_axis_cw_tdata(1 downto 0) /= "10" then
                                       delaylast         <= '1';
                                    elsif s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+2) = '1' and 
                                       s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+3) = '1' then
                                       delaylast         <= '1';
                                    end if;
                                 end if;
                                 if tlppipeline /= "100" then
                                    wrreqsetsig   <= '1';
                                    wrreqpendsig <= wrreqpendsig + 1;
                                    if s_axis_cw_tdata(29) = '0' then
                                       if s_axis_cw_tlast = '1' then
                                          wrreqsmsig       <= onedwlength;
                                          s_axis_cw_treadysig <= '0';
                                       else
                                          wrreqsmsig  <= datatransfer;
                                          dataoffset  <= '1';
                                       end if;
                                    else
                                       wrreqsmsig  <= datatransfer;
                                    end if;
                                    dataen         <= '1';
                                 else
                                    wrreqsmsig       <= throttle;
                                    s_axis_cw_treadysig <= '0';
                                 end if;
                              else
                                 if s_axis_cw_tlast = '0' then
                                    wrreqsmsig       <= zerolenwr;
                                 else
                                    wrreqsmsig    <= memwrreq;
                                 end if;
                              end if;
                           else
                              if s_axis_cw_tlast = '0' then
                                 wrreqsmsig       <= poisoneddataclkout;
                              else
                                 wrreqsmsig    <= memwrreq;
                              end if;
                              master_int    <= '1';
                           end if;
                        --else
                        --   wrreqsmsig       <= memwrreq;
                        end if;
                     --else
                     --   wrreqsmsig          <= memwrreq;
                     end if;
                  end if;
                  blk_lnk_upsig  <= '0';
               end if;

            when zerolenwr =>
               if blk_lnk_up = '1' then
                  -- Nam - enhance core does not throttle
                  -- coverage off -item b 1 -allfalse
                  if s_axis_cw_tvalid = '1' then
                     if s_axis_cw_tlast = '1' then
                        wrreqsmsig       <= memwrreq;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - zero length write while link_down
               -- coverage off
               else
                  if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                     wrreqsmsig       <= memwrreq;
                  else
                     wrreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on

            when onedwlength =>
               wrreqsetsig <= '0';
               if almost_full = '0' then
               if addroffset3 = '0' and addroffset2 = '0' and addroffset1 = '0' then
                  datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= x"0000_0000_0000_0000_0000_0000" & tempdatareg;
               elsif addroffset3 = '0' and addroffset2 = '0' and addroffset1 = '1' then
                  datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= x"0000_0000_0000_0000" & tempdatareg & x"0000_0000";
               elsif addroffset3 = '0' and addroffset2 = '1' and addroffset1 = '0' then
                  datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= x"0000_0000" & tempdatareg & x"0000_0000_0000_0000";
               elsif addroffset3 = '1' and addroffset2 = '0' and addroffset1 = '0' then
                  datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= tempdatareg & x"0000_0000_0000_0000_0000_0000";
               end if;
               datain(C_S_AXIS_DATA_WIDTH)   <= '1';
               wrreqsmsig  <= memwrreq;
               delaylast    <= '0';
               s_axis_cw_treadysig <= '1';
               dataen      <= '0';
               dataoffset  <= '0';
               addroffset1 <= '0';
               addroffset2 <= '0';
               addroffset3 <= '0';
               s_axis_cw_tlasttemp <= s_axis_cw_tlast;
               end if;
            
            when poisoneddataclkout =>
               master_int <= '0';
               if blk_lnk_up = '1' then
                  -- Nam - enhance bridge wont throttle
                  -- coverage off -item b 1 -allfalse
                  if s_axis_cw_tvalid = '1' then
                     if s_axis_cw_tlast = '1' then
                        wrreqsmsig <= memwrreq;
                     end if;
                  end if;
               -- Nam -- extremely hard to hit case - poison data while linkdown
               -- coverage off                  
               else
                  if s_axis_cw_tvalid = '1' and s_axis_cw_tlast = '1' then
                     wrreqsmsig       <= memwrreq;
                  else
                     wrreqsmsig       <= blklinkdown;
                  end if;
               end if;
               -- coverage on
            
            when blklinkdown =>
               -- Nam - enhance bridge wont throttle
               -- coverage off -item b 1 -allfalse            
               if s_axis_cw_tvalid = '1' then
                  if s_axis_cw_tlast = '1' then
                     wrreqsmsig     <= idle;
                  end if;
               -- CR 655336
               -- MWr TLP may finish in single beat so there won't be further valids/last beat
               else
                  wrreqsmsig     <= idle;
               end if;

            when throttle =>
               if blk_lnk_up = '1' then
                  if tlppipeline /= "100" then
                     wrreqsetsig      <= '1';
                     wrreqpendsig <= wrreqpendsig + 1;
                     s_axis_cw_treadysig <= '1';
                     if tlpfmtsig(0) = '0' then
                        if s_axis_cw_tlasttemp = '1' then
                           wrreqsmsig       <= onedwlength;
                           s_axis_cw_treadysig <= '0';
                        else
                           wrreqsmsig       <= datatransfer;
                           dataoffset       <= '1';
                        end if;
                     else
                        wrreqsmsig <= datatransfer;
                     end if;
                     dataen        <= '1';
                  end if;
               -- Nam -- extremely hard to hit case. We covered this with the weekend run - 10 hits
               -- coverage off
               else
                  wrreqsmsig    <= blklinkdown;
                  s_axis_cw_treadysig <= '1';
               end if;
               -- coverage on

            when datatransfer =>
               wrreqsetsig <= '0';
               -- Nam - enhance bridge wont throttle -  -- tool issue, work work when the if statement is more than 1 line
               -- coverage off -item bc 1 -allfalse -condrow 3
               if s_axis_cw_tvalid = '1' or s_axis_cw_tlasttemp = '1' then
                  s_axis_cw_treadysig <= not(almost_full);
                  if almost_full = '0' then
                  if s_axis_cw_treadysig = '1' or s_axis_cw_tlasttemp = '1' then
                  if dataoffset  = '1' then
                     if addroffset1 = '0' and addroffset2 = '0' and addroffset3 = '0' then
                        datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                           little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                             C_S_AXIS_DATA_WIDTH/2)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 
                               C_S_AXIS_DATA_WIDTH/4)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) 
                                    & tempdatareg;
                        tempdatareg <= 
                           little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                             C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4));
                     else
                        if addroffset1 = '1' then
                           if padzeroes = '0' then
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto C_S_AXIS_DATA_WIDTH/4)) & 
                                    little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & 
                                    s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2-1 downto 0);
                           else
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto C_S_AXIS_DATA_WIDTH/4)) & 
                                    little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & 
                                    tempdatareg & x"00000000";
                              padzeroes <= '0';
                           end if;
                           s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2-1 downto 0) <= 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4)) & 
                                  little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                                    C_S_AXIS_DATA_WIDTH/2));
                           end if;
                           if addroffset2 = '1' then
                           if padzeroes = '0' then
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & 
                                    s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 0);
                           else
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & tempdatareg & 
                                   x"0000000000000000";
                              padzeroes <= '0';
                           end if;
                           s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 0) <= 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4)) & 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                                   C_S_AXIS_DATA_WIDTH/2)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 
                                     C_S_AXIS_DATA_WIDTH/4));
                           end if;
                           if addroffset3 = '1' then
                           if padzeroes = '0' then
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= s_axis_cw_tdatatemp;
                           else
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= tempdatareg & x"000000000000000000000000";
                              padzeroes <= '0';
                           end if;
                           s_axis_cw_tdatatemp <= little_to_big_endian32(s_axis_cw_tdata(127 downto 96)) & 
                              little_to_big_endian32(s_axis_cw_tdata(95 downto 64)) & 
                                 little_to_big_endian32(s_axis_cw_tdata(63 downto 32)) & 
                                    little_to_big_endian32(s_axis_cw_tdata(31 downto 0));
                        end if;
                     end if;
                  else
                     if addroffset1 = '0' and addroffset2 = '0' and addroffset3 = '0' then
                        datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= little_to_big_endian32(s_axis_cw_tdata(127 downto 96)) & 
                           little_to_big_endian32(s_axis_cw_tdata(95 downto 64)) & 
                              little_to_big_endian32(s_axis_cw_tdata(63 downto 32)) & 
                                 little_to_big_endian32(s_axis_cw_tdata(31 downto 0));
                     else
                        if addroffset1 = '1' then
                           if padzeroes = '0' then
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                                   C_S_AXIS_DATA_WIDTH/2)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 
                                     C_S_AXIS_DATA_WIDTH/4)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 
                                       downto 0)) & s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/4-1 downto 0);
                           else
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                                   C_S_AXIS_DATA_WIDTH/2)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto 
                                     C_S_AXIS_DATA_WIDTH/4)) & little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 
                                       downto 0)) & x"00000000";
                              padzeroes <= '0';
                           end if;
                           s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/4-1 downto 0) <= 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4));
                        end if;
                        if addroffset2 = '1' then
                           if padzeroes = '0' then
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto C_S_AXIS_DATA_WIDTH/4)) & 
                                    little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & 
                                    s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2-1 downto 0);
                           else
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto C_S_AXIS_DATA_WIDTH/4)) & 
                                    little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & x"0000000000000000";
                              padzeroes <= '0';
                           end if;
                           s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2-1 downto 0) <= 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4)) & 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                                   C_S_AXIS_DATA_WIDTH/2));
                        end if;
                        if addroffset3 = '1' then
                           if padzeroes = '0' then
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & 
                                    s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 0);
                           else
                              datain(C_S_AXIS_DATA_WIDTH-1 downto 0) <= 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/4-1 downto 0)) & 
                                   x"000000000000000000000000";
                              padzeroes <= '0';
                           end if;
                           s_axis_cw_tdatatemp(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 0) <= 
                              little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH-1 downto 
                                C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4)) & 
                                 little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2+C_S_AXIS_DATA_WIDTH/4-1 downto 
                                   C_S_AXIS_DATA_WIDTH/2)) & 
                                    little_to_big_endian32(s_axis_cw_tdata(C_S_AXIS_DATA_WIDTH/2-1 downto C_S_AXIS_DATA_WIDTH/4));
                        end if;
                     end if;
                  end if;
                  if delaylast = '0' then
                     datain(C_S_AXIS_DATA_WIDTH) <= s_axis_cw_tlast;
                     if s_axis_cw_tlast = '1' then
                        wrreqsmsig  <= memwrreq;
                        dataen      <= '0';
                        dataoffset  <= '0';
                        addroffset1 <= '0';
                        addroffset2 <= '0';
                        addroffset3 <= '0';
                     end if;
                  else
                     s_axis_cw_tlasttemp <= s_axis_cw_tlast;
                     datain(C_S_AXIS_DATA_WIDTH) <= s_axis_cw_tlasttemp;
                     if s_axis_cw_tlast = '1' then
                        s_axis_cw_treadysig <= '0';
                     end if;
                     if s_axis_cw_tlasttemp = '1' then
                        s_axis_cw_treadysig <= '1';
                        wrreqsmsig <= memwrreq;
                        s_axis_cw_tlasttemp <= '0';
                        dataen      <= '0';
                        dataoffset  <= '0';
                        addroffset1 <= '0';
                        addroffset2 <= '0';
                        addroffset3 <= '0';
                        delaylast   <= '0';
                     end if;
                  end if;
                  end if;
                  end if;
               end if;
               if blk_lnk_up = '0' then
                  blk_lnk_upsig <= '1';
               end if;

            -- coverage off
            when others =>
               wrreqsmsig <= idle;
            -- coverage on
         end case;
      end if;
   end if;
end process;
end generate;

tlplength          <= tlplengthsig;
firstdwbe          <= firstdwbesig;
lastdwbe           <= lastdwbesig;
wrreqset           <= wrreqsetsig;
treadydataenadjust <= s_axis_cw_tlasttemp;
s_axis_cw_tready   <=
   s_axis_cw_treadysig when almost_full = '0' else
   '0';

wrreqpend <= wrreqpendsig;

end behavioral;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_mm_s_masterbridge_rd.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge read function. 
--                   
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_mm_s_masterbridge_rd.vhd
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library xpm;
use xpm.vcomponents.all;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

--library AMDCoreLib;
--use AMDCoreLib.all;

--library UNISIM;
--use UNISIM.VComponents.all;

entity axi_mm_s_masterbridge_rd is
   generic(
      --Family Generics
      C_FAMILY                : string;
      C_M_AXI_ADDR_WIDTH      : integer;
      C_M_AXI_DATA_WIDTH      : integer;
      C_S_AXIS_DATA_WIDTH     : integer;
      C_PCIEBAR_NUM           : integer;
      C_PCIEBAR_AS            : integer;
      C_PCIEBAR_LEN_0         : integer;
      C_PCIEBAR2AXIBAR_0      : std_logic_vector;
      C_PCIEBAR2AXIBAR_0_SEC  : integer;
      C_PCIEBAR_LEN_1         : integer;
      C_PCIEBAR2AXIBAR_1      : std_logic_vector;
      C_PCIEBAR2AXIBAR_1_SEC  : integer;
      C_PCIEBAR_LEN_2         : integer;
      C_PCIEBAR2AXIBAR_2      : std_logic_vector;
      C_PCIEBAR2AXIBAR_2_SEC  : integer;
      C_S_AXIS_USER_WIDTH     : integer;
      C_TRN_NP_FC             : string
      );
   port(
      --AXI Global
      aclk             : in  std_logic; --meaningful port name
      reset            : in  std_logic; --meaningful port name
      --AXI Master Read Address Channel
      m_axi_araddr     : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      m_axi_arlen      : out std_logic_vector(7 downto 0); --meaningful port name
      m_axi_arsize     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_arburst    : out std_logic_vector(1 downto 0); --meaningful port name
      m_axi_arprot     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_arvalid    : out std_logic; --meaningful port name
      m_axi_arready    : in  std_logic; --meaningful port name
      m_axi_arlock     : out std_logic; --meaningful port name
      m_axi_arcache    : out std_logic_vector(3 downto 0); --meaningful port name
      --AXI Master Read Data Channel
      m_axi_rdata      : in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axi_rresp      : in  std_logic_vector(1 downto 0); --meaningful port name
      m_axi_rlast      : in  std_logic; --meaningful port name
      m_axi_rvalid     : in  std_logic; --meaningful port name
      m_axi_rready     : out std_logic; --meaningful port name
      --AXIS Read Target Channel
      s_axis_cr_tdata  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      s_axis_cr_tstrb  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      s_axis_cr_tlast  : in  std_logic; --meaningful port name
      s_axis_cr_tvalid : in  std_logic; --meaningful port name
      s_axis_cr_tready : out std_logic; --meaningful port name
      s_axis_cr_tuser  : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --AXIS Completion Target Channel
      m_axis_cc_tdata  : out std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axis_cc_tstrb  : out std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      m_axis_cc_tlast  : out std_logic; --meaningful port name
      m_axis_cc_tvalid : out std_logic; --meaningful port name
      m_axis_cc_tready : in  std_logic; --meaningful port name
      m_axis_cc_tuser  : out std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --Master Bridge Interrupt Strobes
      master_int_rd    : out std_logic_vector(1 downto 0); --meaningful port name
      --AXI Streaming Block Interface
      blk_lnk_up          : in  std_logic; --meaningful port name
      blk_lnk_up_latch    : out std_logic; --meaningful port name
      blk_dcontrol        : in  std_logic_vector(15 downto 0); --meaningful port name
      blk_bus_number      : in  std_logic_vector(7 downto 0); --meaningful port name
      blk_device_number   : in  std_logic_vector(4 downto 0); --meaningful port name
      blk_function_number : in  std_logic_vector(2 downto 0); --meaningful port name
      --Internal Interface Ordering
      rdreq               : in  std_logic; --meaningful port name
      rdreq_ordernotreq   : out std_logic; --meaningful port name
      orrdreqpipeline     : in std_logic_vector(2 downto 0); --meaningful port name
      slwrreqpend         : in  std_logic_vector(1 downto 0); --meaningful port name
      rdtargetpipeline    : out std_logic_vector(2 downto 0); --meaningful port name
      rdndreqpipeline     : out std_logic_vector(2 downto 0); -- Used in NP OK mode
      rdreqpipeline       : out std_logic_vector(2 downto 0); -- Used in NP OK mode
      np_pkt_complete     : out std_logic_vector(1 downto 0); -- Used in NP Req mode. bit[1] = rdndreqpipeline; bit[0] = rdreqpipeline
      cplpendcpl          : in  cplpendcpl_array; --meaningful port name
      wrpending           : out wrpend_array; --meaningful port name
      wrreqpend           : in  std_logic_vector(2 downto 0); --meaningful port name
      slwrreqpending      : out slwrreqpending_array; --meaningful port name
      compready           : out std_logic_vector(2 downto 0); --meaningful port name
      wrreqcomp           : in  std_logic_vector(2 downto 0); --meaningful port name
      slv_write_idle      : in  std_logic; --meaningful port name
      s_axi_awvalid       : in  std_logic;
      master_wr_idle      : in  std_logic --meaningful port name
      );
end axi_mm_s_masterbridge_rd;

architecture behavioral of axi_mm_s_masterbridge_rd is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

signal sreset, m_axi_rreadysig  : std_logic;
signal dataensig                : std_logic;
signal emptysig, almost_fullsig : std_logic;
signal dinsig, doutsig          : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
signal rd_ensig, wr_ensig       : std_logic;
signal tlpaddrlsig              : tlpaddrl_array;
signal tlplengthsig             : tlplength_array;
signal rrespsig                 : rresp_array;
signal s_axis_cr_tusersig       : barhit_array;
signal bram_depth               : integer range 256 to 4096;
signal sig_rdtargetpipeline     : std_logic_vector(2 downto 0);
signal sig_addrstreampipeline   : std_logic_vector(2 downto 0);

begin

   comp_read_data_fifo : xpm_fifo_sync
   generic map (
     FIFO_MEMORY_TYPE         => "block",
     ECC_MODE                 => "no_ecc",
     FIFO_WRITE_DEPTH         => 1024*128/C_S_AXIS_DATA_WIDTH,
     WRITE_DATA_WIDTH         => C_S_AXIS_DATA_WIDTH,
     PROG_FULL_THRESH         => 10,
     FULL_RESET_VALUE         => 1,
     READ_MODE                => "fwft",
     FIFO_READ_LATENCY        => 0,
     READ_DATA_WIDTH          => C_S_AXIS_DATA_WIDTH,
     USE_ADV_FEATURES         => "1F1F",
     PROG_EMPTY_THRESH        => 10,
     DOUT_RESET_VALUE         => "0",
     WAKEUP_TIME              => 0
     )
   port map (
     rst              => sreset,
     wr_clk           => aclk,
     wr_en            => wr_ensig,
     wr_ack           => open,
     din              => dinsig,
     full             => open,
     almost_full      => almost_fullsig,
     overflow         => open,
     rd_en            => rd_ensig,
     dout             => doutsig,
     empty            => emptysig,
     almost_empty     => open,
     data_valid       => open,
     underflow        => open,
     wr_data_count    => open,
     sleep            => '0',
     injectsbiterr    => '0',
     injectdbiterr    => '0'
     );



comp_axi_s_masterbridge_rd : entity axi_pcie_v2_9_14.axi_s_masterbridge_rd
   generic map(
      --Family Generics
      C_FAMILY            => C_FAMILY,
      C_S_AXIS_DATA_WIDTH => C_S_AXIS_DATA_WIDTH,
      C_S_AXIS_USER_WIDTH => C_S_AXIS_USER_WIDTH,
      C_PCIEBAR_NUM       => C_PCIEBAR_NUM,
      C_PCIEBAR_AS        => C_PCIEBAR_AS,
      C_TRN_NP_FC         => C_TRN_NP_FC
      )
   port map(
      --AXI Global
      aclk             => aclk,
      reset            => reset,
      --AXIS Read Target Channel
      s_axis_cr_tdata  => s_axis_cr_tdata,
      s_axis_cr_tstrb  => s_axis_cr_tstrb,
      s_axis_cr_tlast  => s_axis_cr_tlast,
      s_axis_cr_tvalid => s_axis_cr_tvalid,
      s_axis_cr_tready => s_axis_cr_tready,
      s_axis_cr_tuser  => s_axis_cr_tuser,
      --AXIS Completion Target Channel
      m_axis_cc_tdata  => m_axis_cc_tdata,
      m_axis_cc_tstrb  => m_axis_cc_tstrb,
      m_axis_cc_tlast  => m_axis_cc_tlast,
      m_axis_cc_tvalid => m_axis_cc_tvalid,
      m_axis_cc_tready => m_axis_cc_tready,
      m_axis_cc_tuser  => m_axis_cc_tuser,
      --AXI Streaming Block Interface
      blk_lnk_up          => blk_lnk_up,
      blk_dcontrol        => blk_dcontrol,
      blk_bus_number      => blk_bus_number,
      blk_device_number   => blk_device_number,
      blk_function_number => blk_function_number,
      --Internal Interface
      rresp           => rrespsig,
      rdreq           => rdreq_ordernotreq,
      empty           => emptysig,
      dout            => doutsig,
      tlpaddrl_out    => tlpaddrlsig,
      tlplength_out   => tlplengthsig,
      rd_en           => rd_ensig,
      --Internal Interface Ordering
      rdtargetpipeline_out => sig_rdtargetpipeline,
      orrdreqpipeline => orrdreqpipeline,
      cplpendcpl      => cplpendcpl,
      wrpending       => wrpending,
      wrreqpend       => wrreqpend,
      slv_write_idle  => slv_write_idle,
      master_wr_idle  => master_wr_idle,
      wrreqcomp       => wrreqcomp,
      addrstreampipeline => sig_addrstreampipeline,
      blk_lnk_up_latch_o => blk_lnk_up_latch,
      rdndreqpipeline_o  => rdndreqpipeline,
      rdreqpipeline_o    => rdreqpipeline,
      np_pkt_complete_o  => np_pkt_complete,
      s_axis_cr_tusersig => s_axis_cr_tusersig
      );

comp_axi_mm_masterbridge_rd : entity axi_pcie_v2_9_14.axi_mm_masterbridge_rd
   generic map(
      --Family Generics
      C_FAMILY             => C_FAMILY,
      C_M_AXI_ADDR_WIDTH      => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH      => C_M_AXI_DATA_WIDTH,
      C_PCIEBAR_NUM           => C_PCIEBAR_NUM,
      C_PCIEBAR_AS            => C_PCIEBAR_AS,
      C_PCIEBAR_LEN_0         => C_PCIEBAR_LEN_0,
      C_PCIEBAR2AXIBAR_0      => C_PCIEBAR2AXIBAR_0,
      C_PCIEBAR2AXIBAR_0_SEC  => C_PCIEBAR2AXIBAR_0_SEC,
      C_PCIEBAR_LEN_1         => C_PCIEBAR_LEN_1,
      C_PCIEBAR2AXIBAR_1      => C_PCIEBAR2AXIBAR_1,
      C_PCIEBAR2AXIBAR_1_SEC  => C_PCIEBAR2AXIBAR_1_SEC,
      C_PCIEBAR_LEN_2         => C_PCIEBAR_LEN_2,
      C_PCIEBAR2AXIBAR_2      => C_PCIEBAR2AXIBAR_2,
      C_PCIEBAR2AXIBAR_2_SEC  => C_PCIEBAR2AXIBAR_2_SEC
      )
   port map(
      --AXI Global
      aclk    => aclk,
      reset   => reset,
      --AXI Master Read Address Channel
      m_axi_araddr     => m_axi_araddr,
      m_axi_arlen      => m_axi_arlen,
      m_axi_arsize     => m_axi_arsize,
      m_axi_arburst    => m_axi_arburst,
      m_axi_arprot     => m_axi_arprot,
      m_axi_arvalid    => m_axi_arvalid,
      m_axi_arready    => m_axi_arready,
      m_axi_arlock     => m_axi_arlock,
      m_axi_arcache    => m_axi_arcache,
      --AXI Master Read Data Channel
      m_axi_rdata      => m_axi_rdata,
      m_axi_rresp      => m_axi_rresp,
      m_axi_rlast      => m_axi_rlast,
      m_axi_rvalid     => m_axi_rvalid,
      m_axi_rready     => m_axi_rreadysig,
      --Master Bridge Interrupt Strobes
      master_int      => master_int_rd,
      --Internal Interface
      rdreq           => rdreq,
      almost_full     => almost_fullsig,
      dataen          => dataensig,
      din             => dinsig,
      tlpaddrl        => tlpaddrlsig,
      tlplength       => tlplengthsig,
      rresp           => rrespsig,
      barhit          => s_axis_cr_tusersig,
      blk_lnk_up      => blk_lnk_up,
      --Internal Interface Ordering
      slwrreqpend     => slwrreqpend,
      slwrreqpending  => slwrreqpending,
      compready       => compready,
      addrstreampipeline => sig_addrstreampipeline,
      s_axi_awvalid   => s_axi_awvalid,
      rdtargetpipeline => sig_rdtargetpipeline,
      master_wr_idle  => master_wr_idle
      );

WriteEnable: process(aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         wr_ensig <= '0';
      else
         wr_ensig <= m_axi_rreadysig and m_axi_rvalid and dataensig;
      end if;
   end if;
end process;

m_axi_rready <= m_axi_rreadysig;
sreset <= not(reset);
rdtargetpipeline <= sig_rdtargetpipeline;

end behavioral;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_mm_s_masterbridge_wr.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge write function. 
--                   
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_mm_s_masterbridge_wr.vhd
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library xpm;
use xpm.vcomponents.all;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;

--library AMDCoreLib;
--use AMDCoreLib.all;

entity axi_mm_s_masterbridge_wr is
   generic(
      --Family Generics
      C_FAMILY                : string;
      C_M_AXI_ADDR_WIDTH      : integer;
      C_M_AXI_DATA_WIDTH      : integer;
      C_S_AXIS_DATA_WIDTH     : integer;
      C_PCIEBAR_NUM           : integer;
      C_PCIEBAR_AS            : integer;
      C_PCIEBAR_LEN_0         : integer;
      C_PCIEBAR2AXIBAR_0      : std_logic_vector;
      C_PCIEBAR2AXIBAR_0_SEC  : integer;
      C_PCIEBAR_LEN_1         : integer;
      C_PCIEBAR2AXIBAR_1      : std_logic_vector;
      C_PCIEBAR2AXIBAR_1_SEC  : integer;
      C_PCIEBAR_LEN_2         : integer;
      C_PCIEBAR2AXIBAR_2      : std_logic_vector;
      C_PCIEBAR2AXIBAR_2_SEC  : integer;
      C_S_AXIS_USER_WIDTH     : integer
      );
   port(
      --AXI Global
      aclk             : in  std_logic; --meaningful port name
      reset            : in  std_logic; --meaningful port name
      --AXI Master Write Address Channel
      m_axi_awaddr     : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      m_axi_awlen      : out std_logic_vector(7 downto 0); --meaningful port name
      m_axi_awsize     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_awburst    : out std_logic_vector(1 downto 0); --meaningful port name
      m_axi_awprot     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_awvalid    : out std_logic; --meaningful port name
      m_axi_awready    : in  std_logic; --meaningful port name
      m_axi_awlock     : out std_logic; --meaningful port name
      m_axi_awcache    : out std_logic_vector(3 downto 0); --meaningful port name
      --AXI Master Write Data Channel
      m_axi_wdata      : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axi_wstrb      : out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0); --meaningful port name
      m_axi_wlast      : out std_logic; --meaningful port name
      m_axi_wvalid     : out std_logic; --meaningful port name
      m_axi_wready     : in  std_logic; --meaningful port name
      --AXI Master Write Response Channel
      m_axi_bresp      : in  std_logic_vector(1 downto 0); --meaningful port name
      m_axi_bvalid     : in  std_logic; --meaningful port name
      m_axi_bready     : out std_logic; --meaningful port name
      --Master Bridge Interrupt Strobes
      master_int_wr    : out std_logic_vector(2 downto 0); --meaningful port name
      --Input from Enhanced PCIe
      blk_lnk_up       : in std_logic; --meaningful port name
      --AXIS Write Target Channel
      s_axis_cw_tdata  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      s_axis_cw_tstrb  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      s_axis_cw_tlast  : in  std_logic; --meaningful port name
      s_axis_cw_tvalid : in  std_logic; --meaningful port name
      s_axis_cw_tready : out std_logic; --meaningful port name
      s_axis_cw_tuser  : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --Internal Interface Ordering
      wrreqpend        : out std_logic_vector(2 downto 0); --meaningful port name
      wrreqcomp        : out std_logic_vector(2 downto 0); --meaningful port name
      master_wr_idle   : out std_logic --meaningful port name
      );
end axi_mm_s_masterbridge_wr;

architecture behavioral of axi_mm_s_masterbridge_wr is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

signal tlplengthsig              : std_logic_vector(9 downto 0);
signal firstdwbesig, lastdwbesig : std_logic_vector(3 downto 0);
signal tlpaddrlsig, tlpaddrhsig  : std_logic_vector(31 downto 0);
signal datainsig                 : std_logic_vector(C_S_AXIS_DATA_WIDTH downto 0);
signal dataoutsig                : std_logic_vector(C_M_AXI_DATA_WIDTH downto 0);
signal wrreqsetsig               : std_logic;
signal rdensig, wrensig          : std_logic;
signal treadydataenadjustsig     : std_logic;
signal emptysig, almost_fullsig  : std_logic;
signal dataensig                 : std_logic;
signal twtreadysig               : std_logic;
signal datacompchecksig          : std_logic;
signal tlppipelinesig            : std_logic_vector(2 downto 0);
signal s_axis_cw_tusersig        : std_logic_vector(C_PCIEBAR_NUM-1 downto 0);
signal sreset                    : std_logic;
signal wrreqpendsig              : std_logic_vector(2 downto 0);
signal wrreqcompsig              : std_logic_vector(2 downto 0);

constant DATA_WIDTH              : std_logic_vector(7 downto 0) := conv_std_logic_vector(C_S_AXIS_DATA_WIDTH, 8);
constant BRAM_DEPTH_MUL_512      : std_logic                    := DATA_WIDTH(6) or DATA_WIDTH(5);
constant BRAM_DEPTH_MULTIPLIER   : std_logic_vector(1 downto 0) := BRAM_DEPTH_MUL_512 & DATA_WIDTH(7);
constant BRAM_DEPTH              : integer range 0 to 512       := conv_integer(BRAM_DEPTH_MULTIPLIER);


begin


comp_write_data_fifo : xpm_fifo_sync
   generic map (
     FIFO_MEMORY_TYPE         => "block",
     ECC_MODE                 => "no_ecc",
     FIFO_WRITE_DEPTH         => 256*BRAM_DEPTH,
     WRITE_DATA_WIDTH         => C_S_AXIS_DATA_WIDTH+1,
     PROG_FULL_THRESH         => 10,
     FULL_RESET_VALUE         => 1,
     READ_MODE                => "fwft",
     FIFO_READ_LATENCY        => 0,
     READ_DATA_WIDTH          => C_S_AXIS_DATA_WIDTH+1,
     USE_ADV_FEATURES         => "1F1F",
     PROG_EMPTY_THRESH        => 10,
     DOUT_RESET_VALUE         => "0",
     WAKEUP_TIME              => 0
     )
   port map (
     rst              => sreset,
     wr_clk           => aclk,
     wr_en            => wrensig,
     wr_ack           => open,
     din              => datainsig,
     full             => open,
     almost_full      => almost_fullsig,
     overflow         => open,
     rd_en            => rdensig,
     dout             => dataoutsig,
     empty            => emptysig,
     almost_empty     => open,
     data_valid       => open,
     underflow        => open,
     wr_data_count    => open,
     sleep            => '0',
     injectsbiterr    => '0',
     injectdbiterr    => '0'
     );

comp_axi_s_masterbridge_wr : entity axi_pcie_v2_9_14.axi_s_masterbridge_wr
   generic map(
      --Family Generics
      C_FAMILY            => C_FAMILY,
      C_S_AXIS_DATA_WIDTH => C_S_AXIS_DATA_WIDTH,
      C_S_AXIS_USER_WIDTH => C_S_AXIS_USER_WIDTH,
      C_PCIEBAR_NUM       => C_PCIEBAR_NUM
      )
   port map(
      --AXI Global
      aclk             => aclk,
      reset            => reset,
      --AXIS Write Target Channel
      s_axis_cw_tdata  => s_axis_cw_tdata,
      s_axis_cw_tstrb  => s_axis_cw_tstrb,
      s_axis_cw_tlast  => s_axis_cw_tlast,
      s_axis_cw_tvalid => s_axis_cw_tvalid,
      s_axis_cw_tready => twtreadysig,
      s_axis_cw_tuser  => s_axis_cw_tuser,
      --Master Bridge Interrupt Strobes
      master_int       => master_int_wr(2),
      --Input from Enhanced PCIe
      blk_lnk_up       => blk_lnk_up,
      --Internal Interface
      tlplength          => tlplengthsig,
      firstdwbe          => firstdwbesig,
      lastdwbe           => lastdwbesig,
      tlpaddrl           => tlpaddrlsig,
      tlpaddrh           => tlpaddrhsig,
      datain             => datainsig,
      wrreqset           => wrreqsetsig,
      datacompcheck      => datacompchecksig,
      tlppipeline        => tlppipelinesig,
      dataen             => dataensig,
      almost_full        => almost_fullsig,
      wrreqpend          => wrreqpendsig,
      treadydataenadjust => treadydataenadjustsig
      );

WriteEnable: process(aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         wrensig <= '0';
      else
         wrensig <= (twtreadysig or (treadydataenadjustsig and not(almost_fullsig))) and 
                    (s_axis_cw_tvalid or treadydataenadjustsig) and dataensig;
      end if;
   end if;
end process;

Bar_Hit: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         s_axis_cw_tusersig <= (others => '0');
      elsif twtreadysig = '1' then
         if C_PCIEBAR_AS = 0 then
            s_axis_cw_tusersig <= s_axis_cw_tuser(C_PCIEBAR_NUM+1 downto 2);
         else
            for i in 0 to C_PCIEBAR_NUM-1 loop
               s_axis_cw_tusersig(i) <= s_axis_cw_tuser(2*(i+1));
            end loop;
         end if;
      end if;
   end if;
end process;

comp_axi_mm_masterbridge_wr : entity axi_pcie_v2_9_14.axi_mm_masterbridge_wr
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_M_AXI_ADDR_WIDTH      => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH      => C_M_AXI_DATA_WIDTH,
      C_PCIEBAR_NUM           => C_PCIEBAR_NUM,
      C_PCIEBAR_AS            => C_PCIEBAR_AS,
      C_PCIEBAR_LEN_0         => C_PCIEBAR_LEN_0,
      C_PCIEBAR2AXIBAR_0      => C_PCIEBAR2AXIBAR_0,
      C_PCIEBAR2AXIBAR_0_SEC  => C_PCIEBAR2AXIBAR_0_SEC,
      C_PCIEBAR_LEN_1         => C_PCIEBAR_LEN_1,
      C_PCIEBAR2AXIBAR_1      => C_PCIEBAR2AXIBAR_1,
      C_PCIEBAR2AXIBAR_1_SEC  => C_PCIEBAR2AXIBAR_1_SEC,
      C_PCIEBAR_LEN_2         => C_PCIEBAR_LEN_2,
      C_PCIEBAR2AXIBAR_2      => C_PCIEBAR2AXIBAR_2,
      C_PCIEBAR2AXIBAR_2_SEC  => C_PCIEBAR2AXIBAR_2_SEC
      )
   port map(
      --AXI Global
      aclk    => aclk,
      reset   => reset,
      --AXI Master Write Address Channel
      m_axi_awaddr    => m_axi_awaddr,
      m_axi_awlen     => m_axi_awlen,
      m_axi_awsize    => m_axi_awsize,
      m_axi_awburst   => m_axi_awburst,
      m_axi_awprot    => m_axi_awprot,
      m_axi_awvalid   => m_axi_awvalid,
      m_axi_awready   => m_axi_awready,
      m_axi_awlock    => m_axi_awlock,
      m_axi_awcache   => m_axi_awcache,
      --AXI Master Write Data Channel
      m_axi_wdata     => m_axi_wdata,
      m_axi_wstrb     => m_axi_wstrb,
      m_axi_wlast     => m_axi_wlast,
      m_axi_wvalid    => m_axi_wvalid,
      m_axi_wready    => m_axi_wready,
      --AXI Master Write Response Channel
      m_axi_bresp     => m_axi_bresp,
      m_axi_bvalid    => m_axi_bvalid,
      m_axi_bready    => m_axi_bready,
      --Master Bridge Interrupt Strobes
      master_int      => master_int_wr(1 downto 0),
      --Internal Interface
      wrreqset        => wrreqsetsig,
      datacompcheck   => datacompchecksig,
      tlplength       => tlplengthsig,
      firstdwbe       => firstdwbesig,
      lastdwbe        => lastdwbesig,
      tlpaddrl        => tlpaddrlsig,
      tlpaddrh        => tlpaddrhsig,
      dout            => dataoutsig,
      rd_en           => rdensig,
      empty           => emptysig,
      tlppipeline     => tlppipelinesig,
      barhit          => s_axis_cw_tusersig(C_PCIEBAR_NUM-1 downto 0),
      --Internal Interface Ordering
      wrreqcomp       => wrreqcompsig
      );

s_axis_cw_tready <= twtreadysig;
sreset <= not(reset);

wrreqpend <= wrreqpendsig;
wrreqcomp <= wrreqcompsig;

master_wr_idle <= '1' when wrreqpendsig = wrreqcompsig else
                  '0';

end behavioral;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_mm_s_masterbridge.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI MM/S master bridge. 
--                   
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_mm_s_masterbridge.vhd
--
-------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_MISC.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

--library AMDCoreLib;
--use AMDCoreLib.all;

--library UNISIM;
--use UNISIM.VComponents.all;

entity axi_mm_s_masterbridge is
   generic(
      --Family Generics
      C_FAMILY                : string := "virtex7";
      C_M_AXI_ADDR_WIDTH      : integer := 32;
      C_M_AXI_DATA_WIDTH      : integer := 32;
      C_S_AXIS_DATA_WIDTH     : integer := 32;
      C_PCIEBAR_NUM           : integer := 3;
      C_PCIEBAR_AS            : integer := 1;
      C_PCIEBAR_LEN_0         : integer := 16;
      C_PCIEBAR2AXIBAR_0      : std_logic_vector := x"70000000";
      C_PCIEBAR2AXIBAR_0_SEC  : integer := 0;
      C_PCIEBAR_LEN_1         : integer := 16;
      C_PCIEBAR2AXIBAR_1      : std_logic_vector := x"80000000";
      C_PCIEBAR2AXIBAR_1_SEC  : integer := 0;
      C_PCIEBAR_LEN_2         : integer := 16;
      C_PCIEBAR2AXIBAR_2      : std_logic_vector := x"80000000";
      C_PCIEBAR2AXIBAR_2_SEC  : integer := 0;
      C_S_AXIS_USER_WIDTH     : integer := 12;
      C_TRN_NP_FC             : string  := "FALSE"
      );
   port(
      --AXI Global
      aclk             : in  std_logic; --meaningful port name
      reset            : in  std_logic; --meaningful port name
      --AXI Master Write Address Channel
      m_axi_awaddr     : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      m_axi_awlen      : out std_logic_vector(7 downto 0); --meaningful port name
      m_axi_awsize     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_awburst    : out std_logic_vector(1 downto 0); --meaningful port name
      m_axi_awprot     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_awvalid    : out std_logic; --meaningful port name
      m_axi_awready    : in  std_logic; --meaningful port name
      m_axi_awlock     : out std_logic; --meaningful port name
      m_axi_awcache    : out std_logic_vector(3 downto 0); --meaningful port name
      --AXI Master Write Data Channel
      m_axi_wdata      : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axi_wstrb      : out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0); --meaningful port name
      m_axi_wlast      : out std_logic; --meaningful port name
      m_axi_wvalid     : out std_logic; --meaningful port name
      m_axi_wready     : in  std_logic; --meaningful port name
      --AXI Master Write Response Channel
      m_axi_bresp      : in  std_logic_vector(1 downto 0); --meaningful port name
      m_axi_bvalid     : in  std_logic; --meaningful port name
      m_axi_bready     : out std_logic; --meaningful port name
      --AXIS Write Target Channel
      s_axis_cw_tdata  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      s_axis_cw_tstrb  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      s_axis_cw_tlast  : in  std_logic; --meaningful port name
      s_axis_cw_tvalid : in  std_logic; --meaningful port name
      s_axis_cw_tready : out std_logic; --meaningful port name
      s_axis_cw_tuser  : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --AXI Master Read Address Channel
      m_axi_araddr     : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0); --meaningful port name
      m_axi_arlen      : out std_logic_vector(7 downto 0); --meaningful port name
      m_axi_arsize     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_arburst    : out std_logic_vector(1 downto 0); --meaningful port name
      m_axi_arprot     : out std_logic_vector(2 downto 0); --meaningful port name
      m_axi_arvalid    : out std_logic; --meaningful port name
      m_axi_arready    : in  std_logic; --meaningful port name
      m_axi_arlock     : out std_logic; --meaningful port name
      m_axi_arcache    : out std_logic_vector(3 downto 0); --meaningful port name
      --AXI Master Read Data Channel
      m_axi_rdata      : in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axi_rresp      : in  std_logic_vector(1 downto 0); --meaningful port name
      m_axi_rlast      : in  std_logic; --meaningful port name
      m_axi_rvalid     : in  std_logic; --meaningful port name
      m_axi_rready     : out std_logic; --meaningful port name
      --AXIS Read Target Channel
      s_axis_cr_tdata  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      s_axis_cr_tstrb  : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      s_axis_cr_tlast  : in  std_logic; --meaningful port name
      s_axis_cr_tvalid : in  std_logic; --meaningful port name
      s_axis_cr_tready : out std_logic; --meaningful port name
      s_axis_cr_tuser  : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --AXIS Completion Target Channel
      m_axis_cc_tdata  : out std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0); --meaningful port name
      m_axis_cc_tstrb  : out std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0); --meaningful port name
      m_axis_cc_tlast  : out std_logic; --meaningful port name
      m_axis_cc_tvalid : out std_logic; --meaningful port name
      m_axis_cc_tready : in  std_logic; --meaningful port name
      m_axis_cc_tuser  : out std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0); --meaningful port name
      --AXI Streaming Block Interface
      blk_lnk_up          : in  std_logic; --meaningful port name
      blk_dcontrol        : in  std_logic_vector(15 downto 0); --meaningful port name
      blk_bus_number      : in  std_logic_vector(7 downto 0); --meaningful port name
      blk_device_number   : in  std_logic_vector(4 downto 0); --meaningful port name
      blk_function_number : in  std_logic_vector(2 downto 0); --meaningful port name
      -- Master Bridge Interrupt Strobes
      MDE_int                 : out std_logic; --meaningful port name
      MSE_int                 : out std_logic; --meaningful port name
      MEP_int                 : out std_logic; --meaningful port name
      --Internal Interface Ordering
      slwrreqpend         : in  std_logic_vector(1 downto 0); --meaningful port name
      slwrreqcomp         : in  std_logic_vector(1 downto 0); --meaningful port name
      wrreqpend           : out std_logic_vector(2 downto 0); --meaningful port name
      wrreqcomp           : out std_logic_vector(2 downto 0); --meaningful port name
      slv_write_idle      : in  std_logic; --meaningful port name
      s_axi_awvalid       : in  std_logic; --meaningful port name
      master_wr_idle      : out std_logic; --meaningful port name
      -- signals used to keep track NP buffer availability
      rdndreqpipeline     : out std_logic_vector(2 downto 0); -- Used in NP OK mode
      rdreqpipeline       : out std_logic_vector(2 downto 0); -- Used in NP OK mode
      np_pkt_complete     : out std_logic_vector(1 downto 0)  -- Used in NP Req mode. bit[1] = rdndreqpipeline; bit[0] = rdreqpipeline
      );
end axi_mm_s_masterbridge;

architecture behavioral of axi_mm_s_masterbridge is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of behavioral : architecture is "yes";

signal rdreq, rdreq_ordernotreq       : std_logic;
signal rdtargetpipeline               : std_logic_vector(2 downto 0);
signal slwrreqpending                 : slwrreqpending_array;
signal compready                      : std_logic_vector(2 downto 0);
signal wrreqpendsig, wrreqcompsig     : std_logic_vector(2 downto 0);
signal orrdreqpipeline, orcplpipeline : std_logic_vector(2 downto 0);
signal cplpendcpl                     : cplpendcpl_array;
signal wrpending                      : wrpend_array;
signal sig_master_wr_idle             : std_logic;
signal master_int_wr                  : std_logic_vector(2 downto 0);
signal master_int_rd                  : std_logic_vector(1 downto 0);
signal blk_lnk_up_latch               : std_logic;
type rdorder_states is (wridle,
                        ordercheckreq);

signal rdorder : rdorder_states;

begin

rd_ordering: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         orrdreqpipeline <= (others => '0');
         rdreq <= '0';
      else
         rdreq <= '0';
         case rdorder is
            when wridle =>
               if sig_master_wr_idle = '1' then
                  rdreq <= rdreq_ordernotreq;
                  rdorder <= wridle;
                  if rdreq_ordernotreq = '1' then
                     orrdreqpipeline <= orrdreqpipeline + 1;
                  end if;
               else
                  rdorder <= ordercheckreq;
               end if;
            
            when ordercheckreq =>
               if rdtargetpipeline /= orrdreqpipeline then
                  if wrpending(conv_integer(orrdreqpipeline(1 downto 0)))(2 downto 0) = wrreqcompsig or 
                    wrpending(conv_integer(orrdreqpipeline(1 downto 0)))(3) = '1' then
                     rdreq <= '1';
                     orrdreqpipeline <= orrdreqpipeline + 1;
                     rdorder <= ordercheckreq;
                  end if;
               elsif sig_master_wr_idle = '1' then
                  rdorder <= wridle;
               end if;
            
            -- coverage off
            when others =>
               rdorder <= wridle;
            -- coverage on
         end case;
         if blk_lnk_up_latch = '0' then
            orrdreqpipeline <= rdtargetpipeline;
            rdreq           <= '0';
         end if;
      end if;
   end if;
end process;

cpl_ordering: process (aclk)
begin
   if rising_edge(aclk) then
      if reset = '0' then
         orcplpipeline <= (others => '0');
         cplpendcpl <= (others => '0');
      else
         if compready /= orcplpipeline then
            cplpendcpl(conv_integer(orcplpipeline(1 downto 0))) <= '0';
            if slwrreqpending(conv_integer(orcplpipeline(1 downto 0))) = slwrreqcomp then
               cplpendcpl(conv_integer(orcplpipeline(1 downto 0))) <= '1';
               orcplpipeline <= orcplpipeline + 1;
            end if;
         end if;
      end if;
      if blk_lnk_up_latch = '0' then
         cplpendcpl <= (others => '0');
      end if;
   end if;
end process;

comp_axi_mm_s_masterbridge_wr: entity axi_pcie_v2_9_14.axi_mm_s_masterbridge_wr
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_M_AXI_ADDR_WIDTH      => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH      => C_M_AXI_DATA_WIDTH,
      C_S_AXIS_DATA_WIDTH     => C_S_AXIS_DATA_WIDTH,
      C_PCIEBAR_NUM           => C_PCIEBAR_NUM,
      C_PCIEBAR_AS            => C_PCIEBAR_AS,
      C_PCIEBAR_LEN_0         => C_PCIEBAR_LEN_0,
      C_PCIEBAR2AXIBAR_0      => C_PCIEBAR2AXIBAR_0,
      C_PCIEBAR2AXIBAR_0_SEC  => C_PCIEBAR2AXIBAR_0_SEC,
      C_PCIEBAR_LEN_1         => C_PCIEBAR_LEN_1,
      C_PCIEBAR2AXIBAR_1      => C_PCIEBAR2AXIBAR_1,
      C_PCIEBAR2AXIBAR_1_SEC  => C_PCIEBAR2AXIBAR_1_SEC,
      C_PCIEBAR_LEN_2         => C_PCIEBAR_LEN_2,
      C_PCIEBAR2AXIBAR_2      => C_PCIEBAR2AXIBAR_2,
      C_PCIEBAR2AXIBAR_2_SEC  => C_PCIEBAR2AXIBAR_2_SEC,
      C_S_AXIS_USER_WIDTH     => C_S_AXIS_USER_WIDTH
      )
   port map(
      --AXI Global
      aclk             => aclk,
      reset            => reset,
      --AXI Master Write Address Channel
      m_axi_awaddr     => m_axi_awaddr,
      m_axi_awlen      => m_axi_awlen,
      m_axi_awsize     => m_axi_awsize,
      m_axi_awburst    => m_axi_awburst,
      m_axi_awprot     => m_axi_awprot,
      m_axi_awvalid    => m_axi_awvalid,
      m_axi_awready    => m_axi_awready,
      m_axi_awlock     => m_axi_awlock,
      m_axi_awcache    => m_axi_awcache,
      --AXI Master Write Data Channel
      m_axi_wdata      => m_axi_wdata,
      m_axi_wstrb      => m_axi_wstrb,
      m_axi_wlast      => m_axi_wlast,
      m_axi_wvalid     => m_axi_wvalid,
      m_axi_wready     => m_axi_wready,
      --AXI Master Write Response Channel
      m_axi_bresp      => m_axi_bresp,
      m_axi_bvalid     => m_axi_bvalid,
      m_axi_bready     => m_axi_bready,
      --Master Bridge Interrupt Strobes
      master_int_wr    => master_int_wr,
      --AXI Streaming Block Interface
      blk_lnk_up       => blk_lnk_up,
      --AXIS Write Target Channel
      s_axis_cw_tdata  => s_axis_cw_tdata,
      s_axis_cw_tstrb  => s_axis_cw_tstrb,
      s_axis_cw_tlast  => s_axis_cw_tlast,
      s_axis_cw_tvalid => s_axis_cw_tvalid,
      s_axis_cw_tready => s_axis_cw_tready,
      s_axis_cw_tuser  => s_axis_cw_tuser,
      --Internal Interface Ordering
      wrreqpend        => wrreqpendsig,
      wrreqcomp        => wrreqcompsig,
      master_wr_idle   => sig_master_wr_idle
      );

comp_axi_mm_s_masterbridge_rd: entity axi_pcie_v2_9_14.axi_mm_s_masterbridge_rd
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_M_AXI_ADDR_WIDTH      => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH      => C_M_AXI_DATA_WIDTH,
      C_S_AXIS_DATA_WIDTH     => C_S_AXIS_DATA_WIDTH,
      C_PCIEBAR_NUM           => C_PCIEBAR_NUM,
      C_PCIEBAR_AS            => C_PCIEBAR_AS,
      C_PCIEBAR_LEN_0         => C_PCIEBAR_LEN_0,
      C_PCIEBAR2AXIBAR_0      => C_PCIEBAR2AXIBAR_0,
      C_PCIEBAR2AXIBAR_0_SEC  => C_PCIEBAR2AXIBAR_0_SEC,
      C_PCIEBAR_LEN_1         => C_PCIEBAR_LEN_1,
      C_PCIEBAR2AXIBAR_1      => C_PCIEBAR2AXIBAR_1,
      C_PCIEBAR2AXIBAR_1_SEC  => C_PCIEBAR2AXIBAR_1_SEC,
      C_PCIEBAR_LEN_2         => C_PCIEBAR_LEN_2,
      C_PCIEBAR2AXIBAR_2      => C_PCIEBAR2AXIBAR_2,
      C_PCIEBAR2AXIBAR_2_SEC  => C_PCIEBAR2AXIBAR_2_SEC,
      C_S_AXIS_USER_WIDTH     => C_S_AXIS_USER_WIDTH,
      C_TRN_NP_FC             => C_TRN_NP_FC
      )
   port map(
      --AXI Global
      aclk             => aclk,
      reset            => reset,
      --AXI Master Read Address Channel
      m_axi_araddr     => m_axi_araddr,
      m_axi_arlen      => m_axi_arlen,
      m_axi_arsize     => m_axi_arsize,
      m_axi_arburst    => m_axi_arburst,
      m_axi_arprot     => m_axi_arprot,
      m_axi_arvalid    => m_axi_arvalid,
      m_axi_arready    => m_axi_arready,
      m_axi_arlock     => m_axi_arlock,
      m_axi_arcache    => m_axi_arcache,
      --AXI Master Read Data Channel
      m_axi_rdata      => m_axi_rdata,
      m_axi_rresp      => m_axi_rresp,
      m_axi_rlast      => m_axi_rlast,
      m_axi_rvalid     => m_axi_rvalid,
      m_axi_rready     => m_axi_rready,
      --Master Bridge Interrupt Strobes
      master_int_rd    => master_int_rd,
      --AXIS Read Target Channel
      s_axis_cr_tdata  => s_axis_cr_tdata,
      s_axis_cr_tstrb  => s_axis_cr_tstrb,
      s_axis_cr_tlast  => s_axis_cr_tlast,
      s_axis_cr_tvalid => s_axis_cr_tvalid,
      s_axis_cr_tready => s_axis_cr_tready,
      s_axis_cr_tuser  => s_axis_cr_tuser,
      --AXIS Completion Target Channel
      m_axis_cc_tdata  => m_axis_cc_tdata,
      m_axis_cc_tstrb  => m_axis_cc_tstrb,
      m_axis_cc_tlast  => m_axis_cc_tlast,
      m_axis_cc_tvalid => m_axis_cc_tvalid,
      m_axis_cc_tready => m_axis_cc_tready,
      m_axis_cc_tuser  => m_axis_cc_tuser,
      --AXI Streaming Block Interface
      blk_lnk_up          => blk_lnk_up,
      blk_lnk_up_latch    => blk_lnk_up_latch,
      blk_dcontrol        => blk_dcontrol,
      blk_bus_number      => blk_bus_number,
      blk_device_number   => blk_device_number,
      blk_function_number => blk_function_number,
      --Internal Interface Ordering
      rdreq            => rdreq,
      rdreq_ordernotreq => rdreq_ordernotreq,
      slwrreqpend      => slwrreqpend,
      rdtargetpipeline => rdtargetpipeline,
      rdndreqpipeline  => rdndreqpipeline,
      rdreqpipeline    => rdreqpipeline,
      np_pkt_complete  => np_pkt_complete,
      orrdreqpipeline  => orrdreqpipeline,
      cplpendcpl       => cplpendcpl,
      wrpending        => wrpending,
      wrreqpend        => wrreqpendsig,
      slwrreqpending   => slwrreqpending,
      compready        => compready,
      wrreqcomp        => wrreqcompsig,
      slv_write_idle   => slv_write_idle,
      s_axi_awvalid    => s_axi_awvalid,
      master_wr_idle   => sig_master_wr_idle
      );

wrreqpend <= wrreqpendsig;
wrreqcomp <= wrreqcompsig;
master_wr_idle   <= sig_master_wr_idle;

MDE_int <= master_int_wr(0) or master_int_rd(0);
MSE_int <= master_int_wr(1) or master_int_rd(1);
MEP_int <= master_int_wr(2);

end behavioral;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        register_block.vhd
--
-- Description:     
--                  
-- This VHDL file is the HDL design file for the AXI slave write bridge. 
--                   
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              register_block.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------

entity register_block is
   generic(
      --Family Generics
      C_FAMILY                : string  :="virtex7";
      C_S_AXI_DATA_WIDTH      : integer := 32;
      C_S_AXI_ADDR_WIDTH      : integer := 32;
      C_AXIBAR_NUM            : integer := 6;
      C_INCLUDE_BAROFFSET_REG : integer := 1;
      C_AXIBAR2PCIEBAR_0       : std_logic_vector:=x"00000000";
      C_AXIBAR2PCIEBAR_1       : std_logic_vector:=x"00000000";
      C_AXIBAR2PCIEBAR_2       : std_logic_vector:=x"00000000";
      C_AXIBAR2PCIEBAR_3       : std_logic_vector:=x"00000000";
      C_AXIBAR2PCIEBAR_4       : std_logic_vector:=x"00000000";
      C_AXIBAR2PCIEBAR_5       : std_logic_vector:=x"00000000";
      C_AXIBAR_AS_0           : integer := 0;
      C_AXIBAR_AS_1           : integer := 0;
      C_AXIBAR_AS_2           : integer := 0;
      C_AXIBAR_AS_3           : integer := 0;
      C_AXIBAR_AS_4           : integer := 0;
      C_AXIBAR_AS_5           : integer := 0
   );
   port(
      -- AXI Global
      s_axi_aclk              : in  std_logic;
      reset                   : in  std_logic;

      -- AXI-Lite Slave IPIC
      IP2Bus_Data             : out std_logic_vector(31 downto 0);
      IP2Bus_WrAck            : out std_logic;
      IP2Bus_RdAck            : out std_logic;
      IP2Bus_Error            : out std_logic;
      Bus2IP_Addr             : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      Bus2IP_Data             : in  std_logic_vector(31 downto 0);
      Bus2IP_RNW              : in  std_logic;
      Bus2IP_BE               : in  std_logic_vector(32/8-1 downto 0);
      Bus2IP_CS               : in  std_logic;
      axibar2pciebar0          : out std_logic_vector(63 downto 0);
      axibar2pciebar1          : out std_logic_vector(63 downto 0);
      axibar2pciebar2          : out std_logic_vector(63 downto 0);
      axibar2pciebar3          : out std_logic_vector(63 downto 0);
      axibar2pciebar4          : out std_logic_vector(63 downto 0);
      axibar2pciebar5          : out std_logic_vector(63 downto 0)
   );
end register_block;

architecture structure of register_block is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

   constant C_VSEC2_CAP         : integer := conv_integer(x"00")/4;
   constant C_VSEC2_HDR         : integer := conv_integer(x"04")/4;
   constant C_AXIBAR2PCIEBAR_0A : integer := conv_integer(x"08")/4;
   constant C_AXIBAR2PCIEBAR_0B : integer := conv_integer(x"0C")/4;
   constant C_AXIBAR2PCIEBAR_1A : integer := conv_integer(x"10")/4;
   constant C_AXIBAR2PCIEBAR_1B : integer := conv_integer(x"14")/4;
   constant C_AXIBAR2PCIEBAR_2A : integer := conv_integer(x"18")/4;
   constant C_AXIBAR2PCIEBAR_2B : integer := conv_integer(x"1C")/4;
   constant C_AXIBAR2PCIEBAR_3A : integer := conv_integer(x"20")/4;
   constant C_AXIBAR2PCIEBAR_3B : integer := conv_integer(x"24")/4;
   constant C_AXIBAR2PCIEBAR_4A : integer := conv_integer(x"28")/4;
   constant C_AXIBAR2PCIEBAR_4B : integer := conv_integer(x"2C")/4;
   constant C_AXIBAR2PCIEBAR_5A : integer := conv_integer(x"30")/4;
   constant C_AXIBAR2PCIEBAR_5B : integer := conv_integer(x"34")/4;

   type axi_bar_array is array (0 to 11) of std_logic_vector(0 to 63);
   type integer_array  is array (0 to 5) of integer range 0 to 1;
   type register_bar_array is array (0 to 11) of std_logic_vector(31 downto 0);

   constant C_AXIBAR_AS_ARRAY : integer_array:=(
      C_AXIBAR_AS_0,
      C_AXIBAR_AS_1,
      C_AXIBAR_AS_2,
      C_AXIBAR_AS_3,
      C_AXIBAR_AS_4,
      C_AXIBAR_AS_5);
   constant C_AXIBAR0_UPPER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_0;
   constant C_AXIBAR0_LOWER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_0;
   constant C_AXIBAR1_UPPER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_1;
   constant C_AXIBAR1_LOWER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_1;
   constant C_AXIBAR2_UPPER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_2;
   constant C_AXIBAR2_LOWER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_2;
   constant C_AXIBAR3_UPPER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_3;
   constant C_AXIBAR3_LOWER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_3;
   constant C_AXIBAR4_UPPER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_4;
   constant C_AXIBAR4_LOWER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_4;
   constant C_AXIBAR5_UPPER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_5;
   constant C_AXIBAR5_LOWER : std_logic_vector(0 to 63):=x"0000000000000000"+C_AXIBAR2PCIEBAR_5;
   constant C_AXIBAR2PCIEBAR_ARRAY : axi_bar_array:=(
      x"0000000000000000"+C_AXIBAR0_UPPER(0 to 31),
      x"0000000000000000"+C_AXIBAR0_LOWER(32 to 63),
      x"0000000000000000"+C_AXIBAR1_UPPER(0 to 31),
      x"0000000000000000"+C_AXIBAR1_LOWER(32 to 63),
      x"0000000000000000"+C_AXIBAR2_UPPER(0 to 31),
      x"0000000000000000"+C_AXIBAR2_LOWER(32 to 63),
      x"0000000000000000"+C_AXIBAR3_UPPER(0 to 31),
      x"0000000000000000"+C_AXIBAR3_LOWER(32 to 63),
      x"0000000000000000"+C_AXIBAR4_UPPER(0 to 31),
      x"0000000000000000"+C_AXIBAR4_LOWER(32 to 63),
      x"0000000000000000"+C_AXIBAR5_UPPER(0 to 31),
      x"0000000000000000"+C_AXIBAR5_LOWER(32 to 63));

   type register_states is (IDLE, REG_ACCESS, WAIT_CS);
   signal register_state : register_states;

   signal sig_axibar2pciebar_array   : axi_bar_array;
   signal sig_axibar2pciebar_reset   : axi_bar_array;
   signal sig_register_bar_array     : register_bar_array;
   constant VSEC2_CAP                : std_logic_vector(31 downto 0) := x"0001_000b";
   constant VSEC2_HDR                : std_logic_vector(31 downto 0) := x"0380_0002";

   signal sig_bus2ip_addr            : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal sig_bus2ip_rnw             : std_logic;
   signal sig_bus2ip_ce              : std_logic_vector(2**4-1 downto 0);
   signal sig_bus2ip_ce_reg          : std_logic_vector(2**4-1 downto 0);
   signal sig_oob                    : std_logic;

begin

   IP2Bus_Error <= '0';

   process(Bus2IP_Addr)
      begin
         sig_bus2ip_ce <= (others => '0');
         sig_bus2ip_ce(conv_integer(Bus2IP_Addr(5 downto 2))) <= '1';
   end process;


    process(s_axi_aclk)
      begin
        if(rising_edge(s_axi_aclk)) then
          if(reset='0') then
            sig_register_bar_array <= (others=> (others => '0'));
            sig_register_bar_array(C_AXIBAR2PCIEBAR_0A-2) <=sig_axibar2pciebar_reset(0)( 0 to 31);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_0B-2) <=sig_axibar2pciebar_reset(0)(32 to 63);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_1A-2) <=sig_axibar2pciebar_reset(1)( 0 to 31);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_1B-2) <=sig_axibar2pciebar_reset(1)(32 to 63);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_2A-2) <=sig_axibar2pciebar_reset(2)( 0 to 31);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_2B-2) <=sig_axibar2pciebar_reset(2)(32 to 63);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_3A-2) <=sig_axibar2pciebar_reset(3)( 0 to 31);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_3B-2) <=sig_axibar2pciebar_reset(3)(32 to 63);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_4A-2) <=sig_axibar2pciebar_reset(4)( 0 to 31);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_4B-2) <=sig_axibar2pciebar_reset(4)(32 to 63);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_5A-2) <=sig_axibar2pciebar_reset(5)( 0 to 31);
            sig_register_bar_array(C_AXIBAR2PCIEBAR_5B-2) <=sig_axibar2pciebar_reset(5)(32 to 63);
            IP2Bus_RdAck               <= '0';
            IP2Bus_WrAck               <= '0';
            IP2Bus_Data                <= (others => '0');
            sig_bus2ip_rnw             <= '0';
            sig_bus2ip_addr            <= (others => '0');
            sig_bus2ip_ce_reg          <= (others => '0');
            sig_oob                    <= '0';
          else
            sig_bus2ip_ce_reg          <= sig_bus2ip_ce;

            IP2Bus_RdAck               <= '0';
            IP2Bus_WrAck               <= '0';
            IP2Bus_Data                <= (others => '0');
            case register_state is
              when IDLE =>
                sig_register_bar_array(0)   <= sig_register_bar_array(0);
		sig_register_bar_array(1)   <= sig_register_bar_array(1);
		if(Bus2IP_CS ='1') then
                   register_state           <= REG_ACCESS;
                   --if(conv_integer(Bus2IP_Addr(12 downto 10))=0) then
                      sig_oob               <= '0';
                   --else
                   --   sig_oob               <= '1';
                   --end if;
                end if;

              when REG_ACCESS =>
                sig_oob   <= sig_oob;
		-- Nam - FALSE branch will not be taken, impossible condition
                -- NAM / JRH Tool bug doesn't exclude the second condition. removed cov off item b 2. Moved cov off.
                -- coverage off -item c 1 -condrow 1 2
                if(bus2ip_CS ='1' and sig_oob='0') then
                    -----------------------------------------------------------------
                    -- Bridge Register Interface Here
                    -----------------------------------------------------------------
                      register_state        <= WAIT_CS;
                      IP2Bus_RdAck          <= Bus2IP_RNW;
                      IP2Bus_WrAck          <= not Bus2IP_RNW;
                      IP2Bus_Data           <= (others => '0');

                      
                      if(C_Include_Baroffset_Reg=1 and Sig_Bus2ip_Ce_Reg(C_VSEC2_CAP)='1') then
                        if(Bus2IP_RNW='0') then
                          null; --read only
                        else
                          Ip2bus_Data <= VSEC2_CAP;
                        end if;
                      end if;
                      if(C_Include_Baroffset_Reg=1 and Sig_Bus2ip_Ce_Reg(C_VSEC2_HDR)='1') then
                        if(Bus2IP_RNW='0') then
                          null; --read only
                        else
                          Ip2bus_Data <= VSEC2_HDR;
                        end if;
                      end if;

                      --translation for bar 0
                      if(C_Include_Baroffset_Reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_0A)='1') then
                        -- Nam - C_AXIBAR_AS_ARRAY(0)=1 will always be TRUE
                        -- coverage off -item c 1 -condrow 2
                        if(Bus2IP_RNW='0' and C_AXIBAR_AS_ARRAY(0)=1) then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_0A-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_0A-2);
                        end if;
                      end if;
                      if(C_Include_Baroffset_Reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_0B)='1') then
                        if(Bus2IP_RNW='0') then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_0B-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_0B-2);
                        end if;
                      end if;

                      --translation for bar 1
                      if(C_Include_Baroffset_Reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_1A)='1' and C_AXIBAR_NUM>1)
                      then
                        if(Bus2IP_RNW='0' and C_AXIBAR_AS_ARRAY(1)=1) then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_1A-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_1A-2);
                        end if;
                      end if;
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_1B)='1' and C_AXIBAR_NUM>1)
                      then
                        if(Bus2IP_RNW='0') then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_1B-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_1B-2);
                        end if;
                      end if;

                      --translation for bar 2
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_2A)='1' and C_AXIBAR_NUM>2)
                      then
                        if(Bus2IP_RNW='0' and C_AXIBAR_AS_ARRAY(2)=1) then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_2A-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_2A-2);
                        end if;
                      end if;
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_2B)='1' and C_AXIBAR_NUM>2)
                      then
                        if(Bus2IP_RNW='0') then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_2B-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_2B-2);
                        end if;
                      end if;

                      --translation for bar 3
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_3A)='1' and C_AXIBAR_NUM>3)
                      then
                        if(Bus2IP_RNW='0' and C_AXIBAR_AS_ARRAY(3)=1) then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_3A-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_3A-2);
                        end if;
                      end if;
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_3B)='1' and C_AXIBAR_NUM>3)
                      then
                        if(Bus2IP_RNW='0') then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_3B-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_3B-2);
                        end if;
                      end if;

                      --translation for bar 4
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_4A)='1' and C_AXIBAR_NUM>4)
                      then
                        if(Bus2IP_RNW='0' and C_AXIBAR_AS_ARRAY(4)=1) then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_4A-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_4A-2);
                        end if;
                      end if;
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_4B)='1' and C_AXIBAR_NUM>4)
                      then
                        if(Bus2IP_RNW='0') then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_4B-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_4B-2);
                        end if;
                      end if;

                      --translation for bar 5
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_5A)='1' and C_AXIBAR_NUM>5)
                      then
                        if(Bus2IP_RNW='0' and C_AXIBAR_AS_ARRAY(5)=1) then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_5A-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_5A-2);
                        end if;
                      end if;
                      if(C_Include_Baroffset_reg=1 and Sig_Bus2ip_Ce_Reg(C_AXIBAR2PCIEBAR_5B)='1' and C_AXIBAR_NUM>5)
                      then
                        if(Bus2IP_RNW='0') then
                          sig_register_bar_array(C_AXIBAR2PCIEBAR_5B-2) <= Bus2IP_Data(31 downto 0);
                        else
                          Ip2bus_Data <=sig_register_bar_array(C_AXIBAR2PCIEBAR_5B-2);
                        end if;
                      end if;

                -- NAM / JRH Tool bug doesn't exclude the second condition. Moved cov off.
                -- coverage off
                else
                  --should only be here if the CS(0) is set and the
                  --address is not within range (aka out of bounds (oob))
                  if(sig_oob = '1') then
                    IP2Bus_WrAck          <= not Bus2IP_RNW;
                    IP2Bus_RdAck          <= Bus2IP_RNW;
                    register_state        <= WAIT_CS;
                  end if;
                  -- coverage on
                end if;
              when WAIT_CS =>
                sig_register_bar_array(0)   <= sig_register_bar_array(0);
		sig_register_bar_array(1)   <= sig_register_bar_array(1);
		sig_oob                  <= sig_oob;
		if(Bus2IP_CS ='0') then
                  register_state        <= IDLE;
                end if;

            end case;
          end if;
        end if;
    end process;


   --AXI to PCIe translation vectors
   -- Crazy looking code to map the generics to the correct registers based on
   -- BAR size (32 or 64bit addresses)
   process(sig_register_bar_array)
   begin
     for i in 0 to 5 loop
       if(i < C_AXIBAR_NUM) then
         if(C_AXIBAR_AS_ARRAY(i)=0) then
           --32bit bar
           sig_axibar2pciebar_array(i)(0  to 31) <= (others => '0');
           sig_axibar2pciebar_array(i)(32 to 63) <= sig_register_bar_array(C_AXIBAR2PCIEBAR_0A-2+i*2+1);
           sig_axibar2pciebar_reset(i)(0  to 31) <= (others => '0');
           sig_axibar2pciebar_reset(i)(32 to 63) <= C_AXIBAR2PCIEBAR_ARRAY(i*2+1)(32 to 63);
         else
           --64bit bar
           sig_axibar2pciebar_array(i)(0  to 31) <= sig_register_bar_array(C_AXIBAR2PCIEBAR_0A-2+i*2);
           sig_axibar2pciebar_array(i)(32 to 63) <= sig_register_bar_array(C_AXIBAR2PCIEBAR_0A-2+i*2+1);
           sig_axibar2pciebar_reset(i)(0  to 31) <= C_AXIBAR2PCIEBAR_ARRAY(i*2)(32 to 63);
           sig_axibar2pciebar_reset(i)(32 to 63) <= C_AXIBAR2PCIEBAR_ARRAY(i*2+1)(32 to 63);
         end if;
       else
         sig_axibar2pciebar_array(i) <= (others => '0');
         sig_axibar2pciebar_reset(i) <= (others => '0');
       end if;
     end loop;
   end process;

   axibar2pciebar0 <= sig_axibar2pciebar_array(0) when C_INCLUDE_BAROFFSET_REG>0
      else x"0000000000000000"+C_AXIBAR2PCIEBAR_0;
   axibar2pciebar1 <= sig_axibar2pciebar_array(1) when C_INCLUDE_BAROFFSET_REG>0
      else x"0000000000000000"+C_AXIBAR2PCIEBAR_1;
   axibar2pciebar2 <= sig_axibar2pciebar_array(2) when C_INCLUDE_BAROFFSET_REG>0
      else x"0000000000000000"+C_AXIBAR2PCIEBAR_2;
   axibar2pciebar3 <= sig_axibar2pciebar_array(3) when C_INCLUDE_BAROFFSET_REG>0
      else x"0000000000000000"+C_AXIBAR2PCIEBAR_3;
   axibar2pciebar4 <= sig_axibar2pciebar_array(4) when C_INCLUDE_BAROFFSET_REG>0
      else x"0000000000000000"+C_AXIBAR2PCIEBAR_4;
   axibar2pciebar5 <= sig_axibar2pciebar_array(5) when C_INCLUDE_BAROFFSET_REG>0
      else x"0000000000000000"+C_AXIBAR2PCIEBAR_5;

end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        slave_read_cpl_tlp.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI slave read bridge. 
--                   
--                  
-- VHDL-Standard:   VHDL'93
--
-------------------------------------------------------------------------------
-- Structure:   
--              slave_read_cpl_tlp.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.conv_std_logic_vector;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

library xpm;
use xpm.vcomponents.all;

entity slave_read_cpl_tlp is
   generic(
      --Family Generics
      C_FAMILY                : string := "virtex7";
      C_AXIREAD_NUM           : integer := 8;
      C_RD_BUFFER_ADDR_SIZE   : integer := 10;
      C_M_AXIS_DATA_WIDTH     : integer := 32
   );
   port(
      -- AXI Global
      aclk                    : in  std_logic;
      reset                   : in  std_logic;

      -- internal interface
      maxreadreqsize          : in  std_logic_vector(2 downto 0);
      m_axis_rr_tlast         : in  std_logic;
      m_axis_rr_tready        : in  std_logic;
      read_req_sent           : in  std_logic;
      tag_sent                : in  std_logic_vector(7 downto 0);
      length_sent             : in  std_logic_vector(9 downto 0);
      rreq_active             : in  std_logic;
      req_active_ptr          : in  integer range 0 to C_AXIREAD_NUM-1;
      data_stream_out         : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      read_data_bram_we       : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      cpl_buffer_addr         : out std_logic_vector(C_RD_BUFFER_ADDR_SIZE-1 downto 0);
      cpl_data_str_done       : out std_logic;
      tag_in_cpl              : out std_logic_vector(7 downto 0);
      tag_cpl_status_clr      : out tag_cpl_status_clr_array;
      req_cpl_pending         : out std_logic;
      cpl_index               : in  integer range 0 to C_AXIREAD_NUM-1;
      rdata_str_done          : in  std_logic;
      rdata_str_start         : in  std_logic;
      first_word_offset       : in  first_word_offset_array;
      unsupported_req         : out std_logic;
      completer_abort         : out std_logic;
      poisoned_req            : out std_logic_vector(C_AXIREAD_NUM-1 downto 0);
      unexpected_cpl          : out std_logic;
      cpl_timer_timeout_strb  : in  std_logic_vector(C_AXIREAD_NUM-1 downto 0);
      rd_req_index_err        : out integer range 0 to C_AXIREAD_NUM-1;
      blk_lnk_up              : in  std_logic;
      header_ep               : in  std_logic;
      reqID                   : in  std_logic_vector(15 downto 0);
      illegal_burst_trns      : in  std_logic;
      bar_error_trns          : in  std_logic;
      total_length_out        : out integer;
      tag_pending_for_cpl     : out std_logic;
      tag_len_active_valid_o  : out std_logic;

      -- AXI Streaming interface
      s_axis_rc_tdata         : in  std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      s_axis_rc_tstrb         : in  std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      s_axis_rc_tlast         : in  std_logic;
      s_axis_rc_tvalid        : in  std_logic;
      s_axis_rc_tready        : out std_logic
   );
end slave_read_cpl_tlp;

   architecture structure of slave_read_cpl_tlp is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

--TLP Header Structure 

-- Fmt  00      Cpl
--      10      CplD
-- Type 01010   always for completion
-- TC   000     always (default)
-- TD   0       always(no digest field)
-- EP   0       data is not poisoned
--      1       data is poisoned
-- Attr 00      always
-- Length       length is inclusive of partial first/last data DWs
-- CplID        Completer ID
-- CS           Completion Status
-- BCM  0       always
-- Byte Count   Remaining bytes to satisfy request
-- ReqID        get from PCIe core block IF
-- Tag          8-bit 
-- Lower Addr   7 lsbs of address for completion

-- CONSTANTS --
   constant STR_DATA_SIZE            : integer := C_M_AXIS_DATA_WIDTH/32;
   constant NUM_STROBES              : integer := C_M_AXIS_DATA_WIDTH/8;
   constant LENGTH_ACTIVE_BRAM_DEPTH : integer := STR_DATA_SIZE*8*C_AXIREAD_NUM;
   constant LENGTH_ACTIVE_BRAM_SIZE  : integer := log2(LENGTH_ACTIVE_BRAM_DEPTH);
   constant CPL_ADDR_COUNT_WIDTH     : integer := log2(STR_DATA_SIZE*256);

   -----------------------------------------------------------------------------
   -- State Machines
   -----------------------------------------------------------------------------

   type rd_cpl_tlpctlSM_STATES is (IDLE,
                                   HEADER_1,
                                   HEADER_2,
                                   HEADER_3,
                                   FIND_TAG_START,
                                   FIND_TAG_WAIT,
                                   CHECK_STATUS,
                                   ERROR,
                                   GET_ERROR_TLP,
                                   LOAD_ADDR_COUNT_1,
                                   LOAD_ADDR_COUNT_2,
                                   FIRST_DATA,
                                   DATA_STR,
                                   DONE_CHECK);
   signal rd_cpl_tlpctlSM_cs      : rd_cpl_tlpctlSM_STATES;
   signal rd_cpl_tlpctlSM_ns      : rd_cpl_tlpctlSM_STATES;

   type rdreq_cpl_correlateSM_STATES is (IDLE,
                                         REQ_ACTIVE,
                                         STROBE);
   signal rdreq_cpl_correlateSM_cs   : rdreq_cpl_correlateSM_STATES;
   signal rdreq_cpl_correlateSM_ns   : rdreq_cpl_correlateSM_STATES;

   -----------------------------------------------------------------------------

   signal fmt                     : std_logic_vector(1 downto 0);
   signal ep                      : std_logic := '0';
   signal length                  : std_logic_vector(9 downto 0);
   signal completer_id            : std_logic_vector(15 downto 0);
   signal cs                      : std_logic_vector(2 downto 0);
   signal byte_count              : std_logic_vector(11 downto 0);
   signal requester_id            : std_logic_vector(15 downto 0);
   signal tag                     : std_logic_vector(7 downto 0) := x"00";
   signal lower_addr              : std_logic_vector(6 downto 0);
   signal tready_int              : std_logic;
   signal header_dw0              : std_logic_vector(31 downto 0);
   signal header_dw0_nxt          : std_logic_vector(31 downto 0);
   signal header_dw1              : std_logic_vector(31 downto 0);
   signal header_dw1_nxt          : std_logic_vector(31 downto 0);
   signal header_dw2              : std_logic_vector(31 downto 0);
   signal header_dw2_nxt          : std_logic_vector(31 downto 0);
   signal first_payload_dw        : std_logic_vector(31 downto 0);
   signal first_payload_dw_nxt    : std_logic_vector(31 downto 0);
   signal tdata_reg               : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
   signal tdata_reg_d             : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
   signal tstrb_reg               : std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
   signal data_str_valid          : std_logic;
   signal last_data_received      : std_logic;
   signal new_data_received       : std_logic;
   signal cpl_data_str_done_int   : std_logic;
   signal cpl_data_str_done_err   : std_logic;


   signal cpl_addr_count          : integer range 0 to 256*STR_DATA_SIZE;
   signal cpl_addr_count_1        : integer range 0 to 256*STR_DATA_SIZE;
   signal cpl_addr_count_nxt      : integer range 0 to 256*STR_DATA_SIZE;
   signal cpl_addr_count_limit    : integer range 0 to 256*STR_DATA_SIZE;
   signal cpl_addr_count_size     : integer range 0 to 8;

   signal cpl_addr_count_en       : std_logic;
   signal cpl_addr_count_done     : std_logic;

   signal cpl_addr_mask           : std_logic_vector(NUM_STROBES/4-1 downto 0);
   signal cpl_addr_mask_nxt       : std_logic_vector(NUM_STROBES/4-1 downto 0);

   signal ic_data_str_mask        : std_logic_vector(NUM_STROBES/4-1 downto 0);
   signal ic_data_str_mask_nxt    : std_logic_vector(NUM_STROBES/4-1 downto 0);

   signal tag_index               : integer range 0 to 31;
   signal tag_index_nxt           : integer range 0 to 31;
   signal tag_index_to            : integer range 0 to 31;
   signal tag_index_sel           : integer range 0 to 31;
   signal rd_req_index            : integer range 0 to C_AXIREAD_NUM-1;
   signal rd_req_index_nxt        : integer range 0 to C_AXIREAD_NUM-1;
   signal rd_req_index_of_to      : integer range 0 to C_AXIREAD_NUM-1;
   signal rd_req_index_sel        : integer range 0 to C_AXIREAD_NUM-1;

   type tag_cpl_status_array is array (0 to C_AXIREAD_NUM-1) of std_logic_vector(0 to 8*STR_DATA_SIZE-1);
   signal tag_cpl_status_int      : tag_cpl_status_clr_array;
   signal tag_cpl_status_at_to    : std_logic_vector(0 to 8*STR_DATA_SIZE-1);
   signal write_strobes           : std_logic_vector(NUM_STROBES-1 downto 0);
   signal cpl_addr_count_inc      : integer range 0 to 4;
   signal extra_write             : integer range 0 to 6;
   signal extra_write_nxt         : integer range 0 to 6;
   signal data_stream_int         : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
--******************************************************************************
   signal cpl_buffer_addr_int     : std_logic_vector(C_RD_BUFFER_ADDR_SIZE-1 downto 0);
--******************************************************************************
   signal maxreadreqsize_adj      : integer range 0 to 5;
   signal tag_match               : std_logic;
   signal tag_match_nxt           : std_logic;
   signal unsupported_req_int     : std_logic;
   signal completer_abort_int     : std_logic;
   signal poisoned_req_nxt        : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal poisoned_req_int        : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal reqID_match             : std_logic;
   signal tag_map_done            : std_logic;
   signal tag_map_start           : std_logic;
   signal tag_len_active_valid    : std_logic;
   signal rr_tready_tvalid_d      : std_logic;
   type tag_array is array (0 to C_AXIREAD_NUM-1, 0 to STR_DATA_SIZE*8-1) of std_logic_vector(9 downto 0);
   type tag_len_index_array is array (0 to C_AXIREAD_NUM-1) of integer range 0 to STR_DATA_SIZE*8;
   signal tag_active              : tag_array;
   signal tag_active_nxt          : tag_array;
   signal tag_len_index           : tag_len_index_array;
   signal tag_len_index_nxt       : tag_len_index_array;
   signal length_active           : std_logic_vector(9 downto 0);
   signal length_active_reg       : std_logic_vector(9 downto 0);
   signal length_active_we        : std_logic_vector(0 downto 0);
   signal length_active_wr_addr   : std_logic_vector(LENGTH_ACTIVE_BRAM_SIZE-1 downto 0);
   signal length_active_rd_addr   : std_logic_vector(LENGTH_ACTIVE_BRAM_SIZE-1 downto 0);
   signal length_active_rd_addr_d : std_logic_vector(LENGTH_ACTIVE_BRAM_SIZE-1 downto 0);
   signal length_active_rd_addr_to : std_logic_vector(LENGTH_ACTIVE_BRAM_SIZE-1 downto 0);
   signal length_active_rd_en     : std_logic;
   signal cpl_addr_count_save     : std_logic_vector(CPL_ADDR_COUNT_WIDTH-1 downto 0);
   signal cpl_addr_count_read     : std_logic_vector(CPL_ADDR_COUNT_WIDTH-1 downto 0);
   signal cpl_addr_count_we       : std_logic_vector(0 downto 0);
   signal cpl_addr_count_rd_en    : std_logic;
   signal cpl_addr_count_rd_en_ord : std_logic;
   signal load_cpl_addr_count     : std_logic;
   signal load_cpl_addr_count_init : std_logic;
   signal cpl_data_str_done_d     : std_logic;
   signal total_length_out_int    : integer;
   signal cpl_length              : std_logic_vector(9 downto 0);
   signal cpl_to_length_sub       : std_logic;
   signal cpl_to_length_sub_rd    : std_logic;
   signal cplsm_idle              : std_logic;
   signal memrdreq_sent           : std_logic;
   signal length_sent_reg         : std_logic_vector(10 downto 0);
   signal cpl_done_without_err    : std_logic;
   signal cpl_timeout_occurred    : std_logic;
   signal cpl_error               : std_logic;

-- This function converts a 32-bit little endian format to big endian format
   function little_to_big_endian32(datain : std_logic_vector(31 downto 0))
         return std_logic_vector is
      variable dataout : std_logic_vector(31 downto 0);
   begin
      dataout := datain(7 downto 0) & datain(15 downto 8) & datain(23 downto 16) & datain(31 downto 24);
      return(dataout);
   end function;

begin

   s_axis_rc_tready      <= tready_int;

   unsupported_req       <= unsupported_req_int;
   completer_abort       <= completer_abort_int;

   cpl_buffer_addr       <= cpl_buffer_addr_int;

   tag_in_cpl            <= tag;
   rd_req_index_err      <= rd_req_index;
   poisoned_req          <= poisoned_req_int;

   tag_len_active_valid_o <= tag_len_active_valid or rr_tready_tvalid_d;

   cpl_data_str_done     <= cpl_data_str_done_int;

   gen_tag_cpl_status_clr_num_rd : for j in 0 to C_AXIREAD_NUM-1 generate
   begin
     gen_tag_cpl_status_clr_str_size_0to32: for k in 0 to STR_DATA_SIZE*8-1 generate
	tag_cpl_status_clr(j)(k) <= '1' when tag_cpl_status_int(j)(k) = '0' else '0';
     end generate;
     gen_str_data_size_2_1: if STR_DATA_SIZE = 2 or STR_DATA_SIZE =1 generate -- added to clear MSB bits in gen1 configuration
     begin
         gen_tag_cpl_status_clr_str_size_msbs0:for k in STR_DATA_SIZE*8 to 31 generate
           tag_cpl_status_clr(j)(k) <= '0';
      	end generate;
     end generate;
   end generate;
  
   clr_in_g2config: if C_AXIREAD_NUM = 4 generate -- added to clear top array in gen2 configuration
     for_j_upperarray: for j in 4 to 7 generate
     for_k_allbits_in_upperarray: for  k in 0 to 31 generate
           tag_cpl_status_clr(j)(k) <= '0';
      end generate;
    end generate;
   end generate;


   maxreadreqsize_adj    <= 3 when STR_DATA_SIZE = 1 and conv_integer(maxreadreqsize) > 3 else
                            4 when STR_DATA_SIZE /= 1 and conv_integer(maxreadreqsize) > 4 else
                            conv_integer(maxreadreqsize);

   cpl_addr_count_size   <= maxreadreqsize_adj + 5 when STR_DATA_SIZE = 1 else
                            maxreadreqsize_adj + 4 when STR_DATA_SIZE = 2 else
                            maxreadreqsize_adj + 3;

   -- Generate the read buffer address for putting completion data into the buffer
   cpl_buffer_addr_int   <= conv_std_logic_vector(rd_req_index, log2(C_AXIREAD_NUM)) &   
                            (SHL(conv_std_logic_vector(tag_index, 8), conv_std_logic_vector(cpl_addr_count_size,4)) +
                            conv_std_logic_vector((cpl_addr_count +
                            first_word_offset(rd_req_index))/STR_DATA_SIZE, 8));

   fmt                   <= header_dw0(30 downto 29);
   cpl_length            <= header_dw0(9 downto 0);
   cs                    <= header_dw1(15 downto 13);
   requester_id          <= header_dw2(31 downto 16);
   tag                   <= header_dw2(15 downto 8);
   lower_addr            <= header_dw2(6 downto 0);
   
   reqID_match           <= '1' when reqID = requester_id else '0';
   
   total_length_out      <= total_length_out_int;

   -- Tally the total length (in DW) of all MemRd TLP requests outstanding and subtract for completions recieved so far
   -- This value is used in the slave_read_req_tlp module fclimit_block logic
   total_length_out_proccess : process(aclk)
   variable no_hit : BOOLEAN;
   begin
      if(rising_edge(aclk)) then
         if(reset = '0' or blk_lnk_up = '0') then
            total_length_out_int        <= 0;
            tag_index_to                <= 0;
            cpl_to_length_sub_rd        <= '0'; 
            cpl_to_length_sub           <= '0'; 
            memrdreq_sent               <= '0';
            cpl_done_without_err        <= '0';
            length_sent_reg             <= (others => '0');
         else
            cpl_to_length_sub           <= cpl_to_length_sub_rd; 
            if cplsm_idle = '1' then
               if (tag_cpl_status_at_to /= (tag_cpl_status_at_to'range => '0')) and cpl_to_length_sub = '0' then
                  no_hit                      := TRUE;
                  for j in 0 to STR_DATA_SIZE*8-1 loop
                     if tag_cpl_status_at_to(j) = '1' and no_hit then
                        no_hit                      := FALSE;
                        tag_index_to                <= j;
                     end if;
                  end loop;
                  cpl_to_length_sub_rd        <= '1'; 
               end if;
            end if;
            if cpl_to_length_sub_rd = '1' then
               cpl_to_length_sub_rd           <= '0';
            end if;
            if cpl_to_length_sub = '1' then
               if tag_active(rd_req_index_of_to, tag_index_to)(9) = '1' or conv_integer(cpl_addr_count_read) = 0 then
                  if length_active = 0 then
                     total_length_out_int        <= total_length_out_int - 1024;
                  else
                     total_length_out_int        <= total_length_out_int - conv_integer(length_active);
                  end if;
               else
                  total_length_out_int        <= total_length_out_int - conv_integer(cpl_addr_count_read);
               end if;
            elsif memrdreq_sent = '1' then
               total_length_out_int        <= total_length_out_int + conv_integer(length_sent_reg);
               memrdreq_sent               <= '0';
            elsif cpl_done_without_err = '1' then
               total_length_out_int        <= total_length_out_int - conv_integer(cpl_length);
               cpl_done_without_err        <= '0';
            end if;
            if tag_len_active_valid = '1' then
               memrdreq_sent               <= '1';
               if length_sent = 0 then
                  length_sent_reg             <= "10000000000";
               else
                  length_sent_reg             <= '0' & length_sent;
               end if;
            end if;
            if cpl_data_str_done_int = '1' and cpl_data_str_done_err = '0' then
               cpl_done_without_err        <= '1';
            end if;
         end if;
      end if;
   end process;

   -- Process the completion TLPs as they are received, detect any error indication and find out if they are expected
   -- and, if so, put the data payload in the correct section of the read data buffer.
   -- Works with the 'sync' process below
   rd_cpl_tlpctlSM_comb : process(rd_cpl_tlpctlSM_cs, header_dw0, header_dw1, header_dw2, first_payload_dw, fmt, cs,
                                  s_axis_rc_tvalid, s_axis_rc_tlast, tdata_reg, tdata_reg_d, last_data_received,
                                  new_data_received, length, tag_index, rd_req_index, cpl_addr_mask, ic_data_str_mask,
                                  tstrb_reg, extra_write, lower_addr, cpl_addr_count, tag_cpl_status_int,tag_active,
                                  tag_match, poisoned_req_int, reqID_match, tag_map_done, cpl_addr_count_read,
                                  length_active_rd_en, tag_cpl_status_at_to)
   begin
      rd_cpl_tlpctlSM_ns          <= rd_cpl_tlpctlSM_cs;
      header_dw0_nxt              <= header_dw0;
      header_dw1_nxt              <= header_dw1;
      header_dw2_nxt              <= header_dw2;
      first_payload_dw_nxt        <= first_payload_dw;
      tready_int                  <= '0';
      data_str_valid              <= '0';
      cpl_data_str_done_int       <= '0';
      cpl_data_str_done_err       <= '0';
      data_stream_int             <= (others => '0');
      write_strobes               <= (others => '1');
      cpl_addr_mask_nxt           <= cpl_addr_mask;
      ic_data_str_mask_nxt        <= ic_data_str_mask;
      cpl_addr_count_en           <= '0';
      cpl_addr_count_inc          <= 1;
      extra_write_nxt             <= 0;
      unsupported_req_int         <= '0';
      completer_abort_int         <= '0';
      unexpected_cpl              <= '0';
      poisoned_req_nxt            <= poisoned_req_int;
      tag_map_start               <= '0';
      load_cpl_addr_count         <= '0';
      load_cpl_addr_count_init    <= '0';
      cpl_addr_count_rd_en        <= '0';
      cplsm_idle                  <= '0';
      cpl_error                   <= '0';
      case rd_cpl_tlpctlSM_cs is
         when IDLE =>
            cplsm_idle            <= '1';
            if (tag_cpl_status_at_to = (tag_cpl_status_at_to'range => '0')) then
               tready_int            <= '1';
            end if;
            if s_axis_rc_tvalid = '1' and (tag_cpl_status_at_to = (tag_cpl_status_at_to'range => '0')) then
               if C_M_AXIS_DATA_WIDTH /= 128 then
                  if s_axis_rc_tlast = '0' then
                     rd_cpl_tlpctlSM_ns    <= HEADER_1;
                  end if;
               else
                  rd_cpl_tlpctlSM_ns    <= HEADER_1;
               end if;
            end if;

         when HEADER_1 =>
            if C_M_AXIS_DATA_WIDTH = 32 then
               header_dw0_nxt        <= tdata_reg;
               tready_int            <= '1';
               if s_axis_rc_tvalid = '1' then
                  if s_axis_rc_tlast = '0' then
                     rd_cpl_tlpctlSM_ns    <= HEADER_2;
                  -- coverage off
                  else
                     rd_cpl_tlpctlSM_ns    <= IDLE;
                  end if;
                  -- coverage on
               end if;
            elsif C_M_AXIS_DATA_WIDTH = 64 then
               header_dw0_nxt        <= tdata_reg(31 downto 0);
               header_dw1_nxt        <= tdata_reg(63 downto 32);
               tready_int            <= '1';
               if s_axis_rc_tvalid = '1' then
                  rd_cpl_tlpctlSM_ns    <= HEADER_2;
               end if;
            else
               header_dw0_nxt        <= tdata_reg(31 downto 0);
               header_dw1_nxt        <= tdata_reg(63 downto 32);
               header_dw2_nxt        <= tdata_reg(95 downto 64);
               first_payload_dw_nxt  <= little_to_big_endian32(tdata_reg(127 downto 96));
               rd_cpl_tlpctlSM_ns    <= FIND_TAG_START;
            end if;

         when HEADER_2 =>
            if C_M_AXIS_DATA_WIDTH = 32 then
               header_dw1_nxt        <= tdata_reg;
               tready_int            <= '1';
               if s_axis_rc_tvalid = '1' then
                  rd_cpl_tlpctlSM_ns    <= HEADER_3;
               end if;
            else
               header_dw2_nxt        <= tdata_reg(31 downto 0);
               first_payload_dw_nxt  <= little_to_big_endian32(tdata_reg(63 downto 32));
               rd_cpl_tlpctlSM_ns    <= FIND_TAG_START;
            end if;

         when HEADER_3 =>
            header_dw2_nxt        <= tdata_reg(31 downto 0);
            rd_cpl_tlpctlSM_ns    <= FIND_TAG_START;

         when FIND_TAG_START =>
            tag_map_start         <= '1';
            if tag_map_done = '1' then
               rd_cpl_tlpctlSM_ns    <= CHECK_STATUS;
            else
               rd_cpl_tlpctlSM_ns    <= FIND_TAG_WAIT;
            end if;

         when FIND_TAG_WAIT =>
            if tag_map_done = '1' then
               rd_cpl_tlpctlSM_ns    <= CHECK_STATUS;
            end if;

         when CHECK_STATUS =>
            if tag_match = '1' and reqID_match = '1' then
               if length_active_rd_en = '1' then 
                  if fmt = "10" and cs = "000" then
                     rd_cpl_tlpctlSM_ns    <= LOAD_ADDR_COUNT_1;
                  else
                     rd_cpl_tlpctlSM_ns    <= ERROR;
                  end if;
               end if;
            else
               unexpected_cpl              <= '1';
               rd_cpl_tlpctlSM_ns          <= GET_ERROR_TLP;
            end if;

         when ERROR =>
            cpl_error                   <= '1';
            if cs = "100" then -- CA status
               completer_abort_int         <= '1';
            elsif cs /= "000" then -- UR status covers reserved as well
               unsupported_req_int         <= '1';
            end if;
            if last_data_received = '0' then
               tready_int                  <= '1';
               rd_cpl_tlpctlSM_ns          <= GET_ERROR_TLP;
            else
               cpl_data_str_done_int       <= '1';
               cpl_data_str_done_err       <= '1';
               rd_cpl_tlpctlSM_ns          <= DONE_CHECK;
            end if;

         when GET_ERROR_TLP => -- clock out remainder of TLP
            cpl_error                   <= '1';
            if last_data_received = '0' then
               tready_int                  <= '1';
            else
               cpl_data_str_done_int       <= '1';
               cpl_data_str_done_err       <= '1';
               rd_cpl_tlpctlSM_ns          <= DONE_CHECK;
            end if;

         when LOAD_ADDR_COUNT_1 =>
            cpl_addr_count_rd_en  <= '1';
            rd_cpl_tlpctlSM_ns    <= LOAD_ADDR_COUNT_2;
         when LOAD_ADDR_COUNT_2 =>
            if C_M_AXIS_DATA_WIDTH = 32 then -- no payload yet for 32-bit
               tready_int            <= '1';
            end if;
            if tag_active(rd_req_index,tag_index)(9) = '1' then
               load_cpl_addr_count_init <= '1';
            else
               load_cpl_addr_count      <= '1';
            end if;
            rd_cpl_tlpctlSM_ns    <= FIRST_DATA;
            if header_dw0(14) = '1' then -- mark request poisoned if ep set
               poisoned_req_nxt(rd_req_index) <= '1';
            end if;
         when FIRST_DATA =>
            data_str_valid        <= '1';
            if C_M_AXIS_DATA_WIDTH = 32 then
               cpl_addr_count_en   <= '1';
               data_stream_int                <= little_to_big_endian32(tdata_reg);
               if last_data_received = '1' then
                  cpl_data_str_done_int <= '1';
                  rd_cpl_tlpctlSM_ns    <= IDLE;
               else
                  tready_int            <= '1';
                  rd_cpl_tlpctlSM_ns    <= DATA_STR;
               end if;
            elsif C_M_AXIS_DATA_WIDTH = 64 then
               cpl_addr_count_en   <= '1';
               ic_data_str_mask_nxt           <= "11";
               if lower_addr(2) = '1' then -- lower address is upper dw
                  write_strobes                  <= x"F0";
                  cpl_addr_mask_nxt   <= "11";
                  data_stream_int                <= first_payload_dw & x"0000_0000";
               else -- new BRAM address 
                  write_strobes                  <= x"0F";
                  cpl_addr_mask_nxt   <= "10"; -- only wrote to lower dw
                  data_stream_int(31 downto 0)   <= first_payload_dw;
               end if;
               if last_data_received = '1' then
                  cpl_data_str_done_int          <= '1';
                  rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
               else
                  tready_int                     <= '1';
                  rd_cpl_tlpctlSM_ns             <= DATA_STR;
               end if;
            else--if C_M_AXIS_DATA_WIDTH = 128 then
               cpl_addr_count_en   <= '1';
               ic_data_str_mask_nxt           <= "1111";
               if lower_addr(3 downto 2) = "01" then -- lower address is dw1
                  write_strobes                  <= x"00F0";
                  cpl_addr_mask_nxt   <= "1100";
                  data_stream_int                <= x"0000_0000_0000_0000" & first_payload_dw & x"0000_0000";
               elsif lower_addr(3 downto 2) = "10" then -- lower address is dw2
                  write_strobes                  <= x"0F00";
                  cpl_addr_mask_nxt   <= "1000";
                  data_stream_int                <= x"0000_0000" & first_payload_dw & x"0000_0000_0000_0000";
               elsif lower_addr(3 downto 2) = "11" then -- lower address is dw3
                  write_strobes                  <= x"F000";
                  cpl_addr_mask_nxt   <= "1111";
                  data_stream_int                <= first_payload_dw & x"0000_0000_0000_0000_0000_0000";
               else -- new BRAM address 
                  write_strobes                  <= x"000F";
                  cpl_addr_mask_nxt   <= "1110"; -- only wrote to lower dw
                  data_stream_int                <= x"0000_0000_0000_0000_0000_0000" & first_payload_dw;
               end if;
               if last_data_received = '1' then
                  cpl_data_str_done_int          <= '1';
                  rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
               else
                  tready_int                     <= '1';
                  rd_cpl_tlpctlSM_ns             <= DATA_STR;
               end if;
            end if;

         when DATA_STR =>
            if last_data_received = '0' then
               tready_int                     <= '1';
            end if;
            if C_M_AXIS_DATA_WIDTH = 32 then
               if new_data_received = '1' then
                  data_stream_int                <= little_to_big_endian32(tdata_reg);
                  data_str_valid                 <= '1';
                  cpl_addr_count_en   <= '1';
                  if last_data_received = '1' then
                     cpl_data_str_done_int          <= '1';
                     rd_cpl_tlpctlSM_ns             <= IDLE;
                  end if;
               end if;
            elsif C_M_AXIS_DATA_WIDTH = 64 then
               if new_data_received = '1' then
                  data_str_valid                 <= '1';
                  cpl_addr_count_en              <= '1';
                  if cpl_addr_mask = "10" then --lower dw at BRAM addr was previously written
                     if ic_data_str_mask = "10" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(63 downto 32)) & x"0000_0000";
                        ic_data_str_mask_nxt           <= "11";
                     else
                        data_stream_int                <= little_to_big_endian32(tdata_reg(31 downto 0)) & x"0000_0000";
                        ic_data_str_mask_nxt           <= "10";
                     end if;
                     write_strobes                  <= x"F0";
                     cpl_addr_mask_nxt   <= "11";
                  else -- new BRAM address 
                     if ic_data_str_mask = "10" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(63 downto 32));
                     else
                        data_stream_int                <= little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0));
                     end if;
                     cpl_addr_count_inc             <= 2;
                  end if;
                  if last_data_received = '1' then
                     if tstrb_reg = x"0F" then -- one dw
                        if ic_data_str_mask = "11" then -- no residual from prior data beat
                           cpl_addr_count_inc             <= 1;
                           if cpl_addr_mask = "10" then
                              write_strobes                  <= x"F0";
                           else
                              write_strobes                  <= x"0F";
                              cpl_addr_mask_nxt   <= "10";
                           end if;
                        else
                           cpl_addr_count_inc             <= 2;
                        end if;
                        cpl_data_str_done_int          <= '1';
                        rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                     else -- two dw received
                        if ic_data_str_mask = "11" and cpl_addr_mask = "11" then
                        -- no residual from prior data beat
                           cpl_data_str_done_int          <= '1';
                           rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                        else
                           extra_write_nxt                <= 1;
                        end if;
                     end if;
                  end if;
               elsif extra_write /= 0 then
                  data_str_valid                 <= '1';
                  data_stream_int                <= x"0000_0000" & little_to_big_endian32(tdata_reg(63 downto 32));
                  write_strobes                  <= x"0F";
                  cpl_addr_count_en   <= '1';
                  ic_data_str_mask_nxt           <= "11";
                  cpl_addr_mask_nxt   <= "10";
                  extra_write_nxt                <= 0;
                  cpl_data_str_done_int          <= '1';
                  rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
               end if;
            else--if C_M_AXIS_DATA_WIDTH = 128 then
               if new_data_received = '1' then
                  data_str_valid                 <= '1';
                  cpl_addr_count_en   <= '1';
                  if cpl_addr_mask = "1110" then --dw0 at BRAM address was previously written
                     if ic_data_str_mask = "1110" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg_d(127 downto 96)) &
                                                          little_to_big_endian32(tdata_reg_d(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg_d(63 downto 32)) & x"0000_0000";
                        ic_data_str_mask_nxt           <= "1111";
                     elsif ic_data_str_mask = "1100" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(127 downto 96)) &
                                                          little_to_big_endian32(tdata_reg_d(95 downto 64)) & x"0000_0000";
                        ic_data_str_mask_nxt           <= "1110";
                     elsif ic_data_str_mask = "1000" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(127 downto 96)) & x"0000_0000";
                        ic_data_str_mask_nxt           <= "1100";
                     else
                        data_stream_int                <= little_to_big_endian32(tdata_reg(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0)) & x"0000_0000";
                        ic_data_str_mask_nxt           <= "1000";
                     end if;
                     cpl_addr_count_inc             <= 3;
                     write_strobes                  <= x"FFF0";
                     cpl_addr_mask_nxt   <= "1111";
                  elsif cpl_addr_mask = "1100" then --dw0, dw1 at BRAM addr were previously written
                     if ic_data_str_mask = "1110" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg_d(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg_d(63 downto 32)) & x"0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1000";
                     elsif ic_data_str_mask = "1100" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg_d(127 downto 96)) &
                                                          little_to_big_endian32(tdata_reg_d(95 downto 64)) & x"0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1111";
                     elsif ic_data_str_mask = "1000" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(127 downto 96)) & x"0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1110";
                     else
                        data_stream_int                <= little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0)) & x"0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1100";
                     end if;
                     cpl_addr_count_inc             <= 2;
                     write_strobes                  <= x"FF00";
                     cpl_addr_mask_nxt   <= "1111";
                  elsif cpl_addr_mask = "1000" then --dw0, dw1, dw2 at BRAM addr were previously written
                     if ic_data_str_mask = "1110" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg_d(63 downto 32)) & x"0000_0000_0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1100";
                     elsif ic_data_str_mask = "1100" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg_d(95 downto 64)) & x"0000_0000_0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1100";
                     elsif ic_data_str_mask = "1000" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg_d(127 downto 96)) & x"0000_0000_0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1111";
                     else
                        data_stream_int                <= little_to_big_endian32(tdata_reg(31 downto 0)) & x"0000_0000_0000_0000_0000_0000";
                        ic_data_str_mask_nxt           <= "1110";
                     end if;
                     write_strobes                  <= x"F000";
                     cpl_addr_mask_nxt   <= "1111";
                  else -- new BRAM addr
                     if ic_data_str_mask = "1110" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(127 downto 96)) &
                                                          little_to_big_endian32(tdata_reg_d(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg_d(63 downto 32));
                        ic_data_str_mask_nxt           <= "1110";
                     elsif ic_data_str_mask = "1100" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(127 downto 96)) &
                                                          little_to_big_endian32(tdata_reg_d(95 downto 64));
                        ic_data_str_mask_nxt           <= "1100";
                     elsif ic_data_str_mask = "1000" then
                        data_stream_int                <= little_to_big_endian32(tdata_reg(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0)) &
                                                          little_to_big_endian32(tdata_reg_d(127 downto 96));
                        ic_data_str_mask_nxt           <= "1000";
                     else
                        data_stream_int                <= little_to_big_endian32(tdata_reg(127 downto 96)) &
                                                          little_to_big_endian32(tdata_reg(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg(63 downto 32)) &
                                                          little_to_big_endian32(tdata_reg(31 downto 0));
                        ic_data_str_mask_nxt           <= "1111";
                     end if;
                     cpl_addr_mask_nxt   <= "1111";
                     cpl_addr_count_inc             <= 4;
                  end if;
                  if last_data_received = '1' then
                     if tstrb_reg = x"000F" then
                        if ic_data_str_mask = "1111" then -- no residual from prior data beat
                           cpl_addr_count_inc             <= 1;
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"000F";
                              cpl_addr_mask_nxt   <= "1110";
                           elsif cpl_addr_mask = "1110" then
                              write_strobes                  <= x"00F0";
                              cpl_addr_mask_nxt   <= "1100";
                           elsif cpl_addr_mask = "1100" then
                              write_strobes                  <= x"0F00";
                              cpl_addr_mask_nxt   <= "1000";
                           else
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                           end if;
                           cpl_data_str_done_int          <= '1';
                           rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                        elsif ic_data_str_mask = "1000" then -- 1 dw of residual data from prior data beat
                           cpl_addr_count_inc             <= 2;
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"00FF";
                              cpl_addr_mask_nxt   <= "1100";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              write_strobes                  <= x"0FF0";
                              cpl_addr_mask_nxt   <= "1000";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1100" then
                              write_strobes                  <= x"FF00";
                              cpl_addr_mask_nxt   <= "1111";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 1;
                           end if;
                        elsif ic_data_str_mask = "1100" then -- 2 dw of residual data from prior data beat
                           cpl_addr_count_inc             <= 3;
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"0FFF";
                              cpl_addr_mask_nxt   <= "1000";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              write_strobes                  <= x"FFF0";
                              cpl_addr_mask_nxt   <= "1111";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 1;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 2;
                           end if;
                        else -- 3 dw of residual data from prior data beat
                           cpl_addr_count_inc             <= 4;
                           cpl_addr_mask_nxt   <= "1111";
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"FFFF";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 2;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 3;
                           end if;
                        end if;
                     elsif tstrb_reg = x"00FF" then
                        if ic_data_str_mask = "1111" then -- no residual from prior data beat
                           cpl_addr_count_inc             <= 2;
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"00FF";
                              cpl_addr_mask_nxt   <= "1100";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              write_strobes                  <= x"0FF0";
                              cpl_addr_mask_nxt   <= "1000";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1100" then
                              write_strobes                  <= x"FF00";
                              cpl_addr_mask_nxt   <= "1111";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 1;
                           end if;
                        elsif ic_data_str_mask = "1000" then -- 1 dw of residual data from prior data beat
                           cpl_addr_count_inc             <= 3;
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"0FFF";
                              cpl_addr_mask_nxt   <= "1000";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              write_strobes                  <= x"FFF0";
                              cpl_addr_mask_nxt   <= "1111";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 1;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 2;
                           end if;
                        elsif ic_data_str_mask = "1100" then -- 2 dw of residual data from prior data beat
                           cpl_addr_count_inc             <= 4;
                           if cpl_addr_mask = "1111" then
                              write_strobes                  <= x"FFFF";
                              cpl_addr_mask_nxt   <= "1111";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 2;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 3;
                           end if;
                        else -- 3 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 2;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 3;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 4;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        end if;
                     elsif tstrb_reg = x"0FFF" then
                        if ic_data_str_mask = "1111" then -- no residual from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"0FFF";
                              cpl_addr_mask_nxt   <= "1000";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              cpl_addr_mask_nxt   <= "1111";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 1;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              cpl_addr_mask_nxt   <= "1111";
                              extra_write_nxt                <= 2;
                           end if;
                        elsif ic_data_str_mask = "1000" then -- 1 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 2;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 3;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        elsif ic_data_str_mask = "1100" then -- 2 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 2;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 3;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 4;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        else -- 3 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              extra_write_nxt                <= 2;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 3;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 4;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 5;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        end if;
                     elsif tstrb_reg = x"FFFF" then
                        if ic_data_str_mask = "1111" then -- no residual from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              cpl_data_str_done_int          <= '1';
                              rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 2;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 3;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        elsif ic_data_str_mask = "1000" then -- 1 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              extra_write_nxt                <= 1;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 2;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 3;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 4;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        elsif ic_data_str_mask = "1100" then -- 2 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              extra_write_nxt                <= 2;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 3;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 4;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 5;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        else -- 3 dw of residual data from prior data beat
                           if cpl_addr_mask = "1111" then
                              cpl_addr_count_inc             <= 4;
                              write_strobes                  <= x"FFFF";
                              extra_write_nxt                <= 3;
                           elsif cpl_addr_mask = "1110" then
                              cpl_addr_count_inc             <= 3;
                              write_strobes                  <= x"FFF0";
                              extra_write_nxt                <= 4;
                           elsif cpl_addr_mask = "1100" then
                              cpl_addr_count_inc             <= 2;
                              write_strobes                  <= x"FF00";
                              extra_write_nxt                <= 5;
                           else
                              cpl_addr_count_inc             <= 1;
                              write_strobes                  <= x"F000";
                              extra_write_nxt                <= 6;
                           end if;
                           cpl_addr_mask_nxt   <= "1111";
                        end if;
                     end if;
                  end if;
               elsif extra_write /= 0 then
                  data_str_valid                 <= '1';
                  cpl_addr_count_en   <= '1';
                  case extra_write is 
                     when 1 =>
                        if ic_data_str_mask = "1000" then
                           data_stream_int                <= x"0000_0000_0000_0000_0000_0000" &
                                                             little_to_big_endian32(tdata_reg(127 downto 96));
                        elsif ic_data_str_mask = "1100" then
                           data_stream_int                <= x"0000_0000_0000_0000_0000_0000" &
                                                             little_to_big_endian32(tdata_reg(95 downto 64));
                        elsif ic_data_str_mask = "1110" then
                           data_stream_int                <= x"0000_0000_0000_0000_0000_0000" &
                                                             little_to_big_endian32(tdata_reg(63 downto 32));
                        end if;
                        cpl_addr_mask_nxt   <= "1110";
                        write_strobes                  <= x"000F";
                        cpl_addr_count_inc             <= 1;
                     when 2 =>
                        if ic_data_str_mask = "1100" then
                           data_stream_int                <= x"0000_0000_0000_0000" &
                                                             little_to_big_endian32(tdata_reg(127 downto 96)) &
                                                             little_to_big_endian32(tdata_reg(95 downto 64));
                        elsif ic_data_str_mask = "1110" then
                           data_stream_int                <= x"0000_0000_0000_0000" &
                                                             little_to_big_endian32(tdata_reg(95 downto 64)) &
                                                             little_to_big_endian32(tdata_reg(63 downto 32));
                        end if;
                        cpl_addr_mask_nxt   <= "1100";
                        write_strobes                  <= x"00FF";
                        cpl_addr_count_inc             <= 2;
                     when 3 =>
                        data_stream_int                <= x"0000_0000" & little_to_big_endian32(tdata_reg(127 downto 96))
                                                          & little_to_big_endian32(tdata_reg(95 downto 64)) &
                                                          little_to_big_endian32(tdata_reg(63 downto 32));
                        cpl_addr_mask_nxt   <= "1100";
                        write_strobes                  <= x"0FFF";
                        cpl_addr_count_inc             <= 3;
                     -- coverage off
                     when others =>
                        null;
                     -- coverage on

                  end case;
                  extra_write_nxt                <= 0;
                  cpl_data_str_done_int          <= '1';
                  rd_cpl_tlpctlSM_ns             <= DONE_CHECK;
               end if;
            end if;

         when DONE_CHECK =>
            rd_cpl_tlpctlSM_ns             <= IDLE;

      end case;
   end process;
      
   -- Process the completion TLPs as they are received, detect any error indication and find out if they are expected
   -- and, if so, put the data payload in the correct section of the read data buffer.
   -- Works with the 'comb' process above
   rd_cpl_tlpctlSM_sync : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            rd_cpl_tlpctlSM_cs    <= IDLE;
            header_dw0            <= (others => '1');
            header_dw1            <= (others => '1');
            header_dw2            <= (others => '1');
            first_payload_dw      <= (others => '0');
            tdata_reg             <= (others => '0');
            tdata_reg_d           <= (others => '0');
            tstrb_reg             <= (others => '0');
            last_data_received    <= '0';
            new_data_received     <= '0';
            cpl_addr_mask         <= (others =>'1');
            ic_data_str_mask      <= (others =>'1');
            extra_write           <= 0;
            poisoned_req_int      <= (others => '0');
         else
            rd_cpl_tlpctlSM_cs    <= rd_cpl_tlpctlSM_ns;
            header_dw0            <= header_dw0_nxt;
            header_dw1            <= header_dw1_nxt;
            header_dw2            <= header_dw2_nxt;
            first_payload_dw      <= first_payload_dw_nxt;
            cpl_addr_mask         <= cpl_addr_mask_nxt;
            ic_data_str_mask      <= ic_data_str_mask_nxt;
            extra_write           <= extra_write_nxt;
            poisoned_req_int      <= poisoned_req_nxt;
            if s_axis_rc_tvalid = '1' and tready_int = '1' then
               for i in 0 to NUM_STROBES-1 loop
                  if s_axis_rc_tstrb(i) = '1' then
                     tdata_reg(i*8+7 downto i*8) <= s_axis_rc_tdata(i*8+7 downto i*8);
                  else
                     tdata_reg(i*8+7 downto i*8) <= (others => '0');
                  end if;
               end loop;
               tdata_reg_d           <= tdata_reg;
               tstrb_reg             <= s_axis_rc_tstrb;
               if s_axis_rc_tlast = '1' then -- and rd_cpl_tlpctlSM_cs /= IDLE then
                  last_data_received    <= '1';
               end if;
               new_data_received     <= '1';
            else
               new_data_received     <= '0';
            end if;
            if cpl_data_str_done_int = '1' then
               last_data_received    <= '0';
            end if;
            if header_ep = '1' then
               poisoned_req_int(cpl_index) <= '0';
            end if;
         end if;
      end if;
   end process;


   data_stream_proc : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            data_stream_out       <= (others => '0');
         else
            data_stream_out       <= data_stream_int;
            if data_str_valid = '1' then
               read_data_bram_we     <= write_strobes;
            else
               read_data_bram_we     <= (others => '0');
            end if;
         end if;
      end if;
   end process;

   -- As MemRd TLPs are generated and sent out, keep track of the tag and length values so that they can be used to
   -- to correlate completion TLPs and tally the amount of data payload needed for each
   rdreq_cpl_correlateSM : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            rdreq_cpl_correlateSM_cs                       <= IDLE;
            tag_active                                     <= (others => (others => (others => '0')));
            tag_len_index                                  <= (others => 0);
            rr_tready_tvalid_d                             <= '0';
         else
            tag_len_active_valid                           <= '0';
            rr_tready_tvalid_d                             <= '0';
            length_active_we                               <= (others => '0');
            case rdreq_cpl_correlateSM_cs is
               when IDLE =>      
                  if rreq_active = '1' and illegal_burst_trns = '0' and bar_error_trns = '0' then
                     rdreq_cpl_correlateSM_cs                       <= REQ_ACTIVE;
                  end if;

               when REQ_ACTIVE =>      
                  if m_axis_rr_tlast = '1' and m_axis_rr_tready = '1' then
                     if tag_len_index(req_active_ptr) < STR_DATA_SIZE*8 then
                        tag_active(req_active_ptr, tag_len_index(req_active_ptr))       <= "11" & tag_sent;
                        length_active_we                               <= (others => '1');
                     end if;
                     rdreq_cpl_correlateSM_cs                       <= STROBE;
                     rr_tready_tvalid_d                             <= '1';
                  end if;

               when STROBE =>      
                  -- pass tag_len_active array entry to completion proccessing
                  tag_len_index(req_active_ptr)                  <= tag_len_index(req_active_ptr) + 1;
                  tag_len_active_valid                           <= '1';
                  if read_req_sent = '1' then
                     rdreq_cpl_correlateSM_cs                       <= IDLE;
                  else
                     rdreq_cpl_correlateSM_cs                       <= REQ_ACTIVE;
                  end if;

            end case;
            if rdata_str_start = '1' then
               if cpl_error = '0' then
                  for i in 0 to STR_DATA_SIZE*8-1 loop
                     tag_active(cpl_index, i)                       <= (others => '0');
                  end loop;
               end if;
               tag_len_index(cpl_index)                       <= 0;
            end if;
            if load_cpl_addr_count_init = '1' then
               tag_active(rd_req_index,tag_index)(9)          <= '0';
            end if;
            -- If full completion count clear active tag entry
            if cpl_addr_count_done = '1' then
               tag_active(rd_req_index, tag_index)        <= (others => '0');
            end if;
            -- If Errors clear active tag entry
            if cpl_to_length_sub = '1' then
               tag_active(rd_req_index_of_to, tag_index_to)  <= (others => '0');
            end if;
         end if;
      end if;
   end process;

   validate_tag : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            tag_pending_for_cpl <= '0';
         else
            tag_pending_for_cpl <= '0';
            for i in 0 to C_AXIREAD_NUM-1 loop
               for j in 0 to STR_DATA_SIZE*8-1 loop
                  if(tag_active(i,j)(9 downto 8) /= "00" and tag_active(i,j)(7 downto 0) = tag_sent) then
                     tag_pending_for_cpl <= '1';
                  end if;
               end loop;
            end loop;
         end if;
      end if;
   end process;

   -- Used to find a tag within the tag_active structure and return rd_req_index and tag_index
   -- Works with 'sync' process below
   cpl_tag_mapping_process : process(tag_map_start, tag_active, tag, rd_req_index, tag_index, tag_match)
   variable match : boolean;
   begin
      rd_req_index_nxt      <= rd_req_index;
      tag_index_nxt         <= tag_index;
      tag_match_nxt         <= tag_match;
      tag_map_done          <= '0';
      if C_AXIREAD_NUM = 8 then
         case rd_req_index is
            when 0 =>
               if tag_map_start = '1' then
                  match                 := FALSE;
                  for i in 0 to STR_DATA_SIZE*8-1 loop
                     if ('1' & tag) = tag_active(0,i)(8 downto 0) then
                        tag_index_nxt         <= i;
                        match                 := TRUE;
                     end if;
                  end loop;
                  if match then
                     tag_map_done          <= '1';
                     tag_match_nxt         <= '1';
                  else
                     rd_req_index_nxt      <= 1;
                  end if;
               end if;
            when 1 to 6 =>
               match                 := FALSE;
               for i in 0 to STR_DATA_SIZE*8-1 loop
                  if ('1' & tag) = tag_active(rd_req_index,i)(8 downto 0) then
                     tag_index_nxt         <= i;
                     match                 := TRUE;
                  end if;
               end loop;
               if match then
                  tag_map_done          <= '1';
                  tag_match_nxt         <= '1';
               else
                  rd_req_index_nxt      <= rd_req_index + 1;
               end if;

            when 7 =>
               match                 := FALSE;
               for i in 0 to STR_DATA_SIZE*8-1 loop
                  if ('1' & tag) = tag_active(rd_req_index,i)(8 downto 0) then
                     tag_index_nxt         <= i;
                     match                 := TRUE;
                  end if;
               end loop;
               if match then
                  tag_match_nxt         <= '1';
               else
                  rd_req_index_nxt      <= 0;
               end if;
               tag_map_done          <= '1';

            -- coverage off
            when others =>
               null;
            -- coverage on

         end case;
      else
         case rd_req_index is
            when 0 =>
               if tag_map_start = '1' then
                  match                 := FALSE;
                  for i in 0 to STR_DATA_SIZE*8-1 loop
                     if ('1' & tag) = tag_active(0,i)(8 downto 0) then
                        tag_index_nxt         <= i;
                        match                 := TRUE;
                     end if;
                  end loop;
                  if match then
                     tag_map_done          <= '1';
                     tag_match_nxt         <= '1';
                  else
                     rd_req_index_nxt      <= 1;
                  end if;
               end if;
            when 1 to 2 =>
               match                 := FALSE;
               for i in 0 to STR_DATA_SIZE*8-1 loop
                  if ('1' & tag) = tag_active(rd_req_index,i)(8 downto 0) then
                     tag_index_nxt         <= i;
                     match                 := TRUE;
                  end if;
               end loop;
               if match then
                  tag_map_done          <= '1';
                  tag_match_nxt         <= '1';
               else
                  rd_req_index_nxt      <= rd_req_index + 1;
               end if;

            when 3 =>
               match                 := FALSE;
               for i in 0 to STR_DATA_SIZE*8-1 loop
                  if ('1' & tag) = tag_active(rd_req_index,i)(8 downto 0) then
                     tag_index_nxt         <= i;
                     match                 := TRUE;
                  end if;
               end loop;
               if match then
                  tag_match_nxt         <= '1';
               else
                  rd_req_index_nxt      <= 0;
               end if;
               tag_map_done          <= '1';

            -- coverage off
            when others =>
               null;
            -- coverage on

         end case;
      end if;
   end process;

   -- Used to find a tag within the tag_active structure and return rd_req_index and tag_index
   -- Works with 'comb' process above
   cpl_tag_mapping_process_sync : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0' or cpl_data_str_done_d = '1') then
            rd_req_index          <= 0;
            tag_index             <= 0;
            tag_match             <= '0';
         else
            rd_req_index          <= rd_req_index_nxt;
            tag_index             <= tag_index_nxt;
            tag_match             <= tag_match_nxt;
         end if;
      end if;
   end process;


   -- Maintain the tag_cpl_status structure to know which MemRd TLPs/tags are pending
   tally_tag_cpl_process : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0' or blk_lnk_up = '0') then
            tag_cpl_status_int          <= (others => (others => '0'));
            tag_cpl_status_at_to        <= (others => '0');
            cpl_timeout_occurred        <= '0';
         elsif tag_len_active_valid = '1' then
            for i in 0 to STR_DATA_SIZE*8-1 loop
               if i = tag_len_index(req_active_ptr) - 1  then
                  tag_cpl_status_int(req_active_ptr)(i) <= '1';
               end if;
            end loop;
         end if;
         if cpl_addr_count_done = '1' then
            tag_cpl_status_int(rd_req_index)(tag_index)   <= '0';
         end if;
         -- Errors that must return arbitrary data to AXI MM have status and counters cleared
         if unsupported_req_int = '1' or completer_abort_int = '1' then
            tag_cpl_status_int(rd_req_index)(tag_index)   <= '0';
            -- capture info for fc count adjust
            if STR_DATA_SIZE = 1 then  -- 32-bit
               tag_cpl_status_at_to        <= SHR(x"80", conv_std_logic_vector(tag_index, 5));
            elsif STR_DATA_SIZE = 2 then -- 64-bit
               tag_cpl_status_at_to        <= SHR(x"8000", conv_std_logic_vector(tag_index, 5));
            else -- 128-bit
               tag_cpl_status_at_to        <= SHR(x"80000000",conv_std_logic_vector(tag_index, 5));
            end if;
            rd_req_index_of_to          <= rd_req_index;
         end if;
         -- Check for completion timer timeouts and clear status and counters
         for j in 0 to C_AXIREAD_NUM-1 loop
            if cpl_timer_timeout_strb(j) = '1' then
               cpl_timeout_occurred        <= '1';
               -- capture info for fc count adjust
               tag_cpl_status_at_to        <= tag_cpl_status_int(j)(0 to 8*STR_DATA_SIZE-1);
               rd_req_index_of_to          <= j;
            end if;
         end loop;
         if cpl_to_length_sub = '1' then
            tag_cpl_status_at_to(tag_index_to) <= '0';
         end if;
         if cpl_timeout_occurred = '1' and (tag_cpl_status_at_to = (tag_cpl_status_at_to'range => '0')) then
            tag_cpl_status_int(rd_req_index_of_to) <= (others => '0');
            cpl_timeout_occurred        <= '0';
         end if;
      end if;
   end process;


   -- Completion address counter. The count value for each tag is saved away to and retrieved from the
   -- cpl_addr_count_bram, as needed, to count down the total length of the MemRd TLP/tag
   cpl_addr_count_limit              <= conv_integer(length_active_reg)
                                        when length_active_reg /= "0000000000"
                                        else 256*STR_DATA_SIZE;
   
   cpl_addr_counter_comb1 : process(cpl_addr_count_1, cpl_addr_count_en, cpl_addr_count_limit, rd_req_index,
                                    tag_index, cpl_addr_count_inc, unsupported_req_int, completer_abort_int,
                                    cpl_timer_timeout_strb, load_cpl_addr_count, load_cpl_addr_count_init,
                                    cpl_addr_count_read)
   begin
      cpl_addr_count_nxt          <= cpl_addr_count_1;
      cpl_addr_count_done         <= '0';
      if load_cpl_addr_count_init = '1' then
         cpl_addr_count_nxt          <= cpl_addr_count_limit;
      elsif load_cpl_addr_count = '1' then
         cpl_addr_count_nxt          <= conv_integer(cpl_addr_count_read);
      end if;
      if cpl_addr_count_en = '1' then
         if cpl_addr_count_1 >= cpl_addr_count_inc then
            if (cpl_addr_count_1 = cpl_addr_count_inc) then
               cpl_addr_count_done         <= '1';
            end if;
            cpl_addr_count_nxt          <= cpl_addr_count_1 - cpl_addr_count_inc;
         end if;
      end if;
      if unsupported_req_int = '1' or completer_abort_int = '1' then
         cpl_addr_count_nxt          <= 0;
      end if;
   end process;

   cpl_addr_counter_sync : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            cpl_addr_count_1         <= 0;
            cpl_addr_count           <= 0;
            cpl_data_str_done_d      <= '0';
            length_active_rd_addr_d  <= (others => '0');
            length_active_reg        <= (others => '0');
         else
            cpl_addr_count_1         <= cpl_addr_count_nxt;
            if cpl_addr_count_1 <= cpl_addr_count_limit then
               cpl_addr_count           <= cpl_addr_count_limit - cpl_addr_count_1;
            end if;
            cpl_data_str_done_d      <= cpl_data_str_done_int;
            length_active_rd_addr_d  <= length_active_rd_addr;
            length_active_reg        <= length_active;
         end if;
      end if;
   end process;


   length_active_wr_addr <= conv_std_logic_vector(req_active_ptr, 3) & conv_std_logic_vector(tag_len_index(req_active_ptr), log2(STR_DATA_SIZE*8))
                               when C_AXIREAD_NUM = 8 else
                               conv_std_logic_vector(req_active_ptr, 2) & conv_std_logic_vector(tag_len_index(req_active_ptr), log2(STR_DATA_SIZE*8));

   rd_req_index_sel <= rd_req_index_of_to when (tag_cpl_status_at_to /= (tag_cpl_status_at_to'range => '0')) and cplsm_idle = '1' else rd_req_index;

   tag_index_sel <= tag_index_to when (tag_cpl_status_at_to /= (tag_cpl_status_at_to'range => '0')) and cplsm_idle = '1' else tag_index;

   length_active_rd_addr <= conv_std_logic_vector(rd_req_index_sel, 3) & conv_std_logic_vector(tag_index_sel, log2(STR_DATA_SIZE*8))
                               when C_AXIREAD_NUM = 8 else
                               conv_std_logic_vector(rd_req_index_sel, 2) & conv_std_logic_vector(tag_index_sel, log2(STR_DATA_SIZE*8));

   length_active_rd_en   <= '0' when length_active_we = "1" else '1';


   comp_length_active_bram : xpm_memory_tdpram
   generic map (
      MEMORY_SIZE        => (LENGTH_ACTIVE_BRAM_DEPTH * 10),
      MEMORY_PRIMITIVE   => "block",               --string; "auto", "distributed", "block" or "ultra" ;
      CLOCKING_MODE      => "common_clock",
      MEMORY_INIT_FILE   => "none",
      MEMORY_INIT_PARAM  => "",
      USE_MEM_INIT       => 1,
      WAKEUP_TIME        => "disable_sleep",
      MESSAGE_CONTROL    => 0,
      ECC_MODE           => "no_ecc",
      AUTO_SLEEP_TIME    => 0,
      -- Port A module generics
      WRITE_DATA_WIDTH_A => 10,
      READ_DATA_WIDTH_A  => 10,
      BYTE_WRITE_WIDTH_A => 10,
      ADDR_WIDTH_A       => LENGTH_ACTIVE_BRAM_SIZE,
      READ_RESET_VALUE_A => "0",
      READ_LATENCY_A     => 1,
      WRITE_MODE_A       => "write_first",
      -- Port B module generics
      WRITE_DATA_WIDTH_B => 10,
      READ_DATA_WIDTH_B  => 10,
      BYTE_WRITE_WIDTH_B => 10,
      ADDR_WIDTH_B       => LENGTH_ACTIVE_BRAM_SIZE,
      READ_RESET_VALUE_B => "0",
      READ_LATENCY_B     => 1,
      WRITE_MODE_B       => "write_first"
      )
   port map (
      sleep          => '0',
      -- Port A module ports
      clka           => aclk,
      rsta           => '0',   
      ena            => length_active_we(0),
      regcea         => '1',
      wea            => length_active_we,
      addra          => length_active_wr_addr,
      dina           => length_sent,
      injectsbiterra => '0',
      injectdbiterra => '0',
      douta          => open,
      sbiterra       => open,
      dbiterra       => open,
      -- Port B module ports
      clkb           => aclk,
      rstb           => '0',  
      enb            => length_active_rd_en,
      regceb         => '1',
      web            => (OTHERS => '0'),
      addrb          => length_active_rd_addr,
      dinb           => (OTHERS => '0'),
      injectsbiterrb => '0',
      injectdbiterrb => '0',
      doutb          => length_active,
      sbiterrb       => open,
      dbiterrb       => open
      );

   cpl_addr_count_save         <= conv_std_logic_vector(cpl_addr_count_1, CPL_ADDR_COUNT_WIDTH);
   cpl_addr_count_we           <= (others => '1') when cpl_done_without_err = '1' and tag_match = '1' else (others => '0');
   cpl_addr_count_rd_en_ord    <= '1' when (tag_cpl_status_at_to /= (tag_cpl_status_at_to'range => '0')) else cpl_addr_count_rd_en; 

   comp_cpl_addr_count_bram : xpm_memory_tdpram
   generic map (
      MEMORY_SIZE        => (LENGTH_ACTIVE_BRAM_DEPTH * CPL_ADDR_COUNT_WIDTH),
      MEMORY_PRIMITIVE   => "block",               --string; "auto", "distributed", "block" or "ultra" ;
      CLOCKING_MODE      => "common_clock",
      MEMORY_INIT_FILE   => "none",
      MEMORY_INIT_PARAM  => "",
      USE_MEM_INIT       => 1,
      WAKEUP_TIME        => "disable_sleep",
      MESSAGE_CONTROL    => 0,
      ECC_MODE           => "no_ecc",
      AUTO_SLEEP_TIME    => 0,
      -- Port A module generics
      WRITE_DATA_WIDTH_A => CPL_ADDR_COUNT_WIDTH,
      READ_DATA_WIDTH_A  => CPL_ADDR_COUNT_WIDTH,
      BYTE_WRITE_WIDTH_A => CPL_ADDR_COUNT_WIDTH,
      ADDR_WIDTH_A       => LENGTH_ACTIVE_BRAM_SIZE,
      READ_RESET_VALUE_A => "0",
      READ_LATENCY_A     => 1,
      WRITE_MODE_A       => "write_first",
      -- Port B module generics
      WRITE_DATA_WIDTH_B => CPL_ADDR_COUNT_WIDTH,
      READ_DATA_WIDTH_B  => CPL_ADDR_COUNT_WIDTH,
      BYTE_WRITE_WIDTH_B => CPL_ADDR_COUNT_WIDTH,
      ADDR_WIDTH_B       => LENGTH_ACTIVE_BRAM_SIZE,
      READ_RESET_VALUE_B => "0",
      READ_LATENCY_B     => 1,
      WRITE_MODE_B       => "write_first"
      )
   port map (
      sleep          => '0',
      -- Port A module ports
      clka           => aclk,
      rsta           => '0',   
      ena            => '1',
      regcea         => '1',
      wea            => cpl_addr_count_we,
      addra          => length_active_rd_addr_d,
      dina           => cpl_addr_count_save,
      injectsbiterra => '0',
      injectdbiterra => '0',
      douta          => open,
      sbiterra       => open,
      dbiterra       => open,
      -- Port B module ports
      clkb           => aclk,
      rstb           => '0',  
      enb            => cpl_addr_count_rd_en_ord,
      regceb         => '1',
      web            => (OTHERS => '0'),
      addrb          => length_active_rd_addr,
      dinb           => (OTHERS => '0'),
      injectsbiterrb => '0',
      injectdbiterrb => '0',
      doutb          => cpl_addr_count_read,
      sbiterrb       => open,
      dbiterrb       => open
      );

end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        slave_read_req_tlp.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI slave read bridge. 
--                   
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              slave_read_req_tlp.vhd
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.conv_std_logic_vector;

--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------



entity slave_read_req_tlp is
   generic(
      --Family Generics
      C_FAMILY                : string  :="virtex7";
      C_S_AXI_ID_WIDTH        : integer := 4;
      C_S_AXI_ADDR_WIDTH      : integer := 32;
      C_S_AXI_DATA_WIDTH      : integer := 32;
      C_M_AXIS_DATA_WIDTH     : integer := 32;
      C_AXIBAR_NUM            : integer := 6;
      C_AXIBAR_0              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0     : std_logic_vector := x"0000_0000";
      C_AXIBAR_1              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1     : std_logic_vector := x"0000_0000";
      C_AXIBAR_2              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2     : std_logic_vector := x"0000_0000";
      C_AXIBAR_3              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3     : std_logic_vector := x"0000_0000";
      C_AXIBAR_4              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4     : std_logic_vector := x"0000_0000";
      C_AXIBAR_5              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5     : std_logic_vector := x"0000_0000";
      C_AXIBAR_AS_0           : integer := 0;
      C_AXIBAR_AS_1           : integer := 0;
      C_AXIBAR_AS_2           : integer := 0;
      C_AXIBAR_AS_3           : integer := 0;
      C_AXIBAR_AS_4           : integer := 0;
      C_AXIBAR_AS_5           : integer := 0;
      C_EP_LINK_PARTNER_RCB   : integer := 0
   );
   port(
      -- AXI Global
      aclk                    : in  std_logic;
      reset                   : in  std_logic;

      -- internal interface
      maxreadreqsize          : in  std_logic_vector(2 downto 0);
      raddr                   : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      length_bytes            : in  std_logic_vector(12 downto 0);
      rbarhit                 : in  std_logic_vector(C_AXIBAR_NUM-1 downto 0);
      araddr_2lsbs            : in  std_logic_vector(1 downto 0);
      last_BE                 : in  std_logic_vector(3 downto 0);
      reqID                   : in  std_logic_vector(15 downto 0);
      req_active              : in  std_logic;
      read_req_sent           : out std_logic;
      tag_sent                : out std_logic_vector(7 downto 0);
      length_sent             : out std_logic_vector(9 downto 0);
      illegal_burst           : in  std_logic;
      illegal_burst_trns      : out std_logic;
      bar_error               : in  std_logic;
      bar_error_trns          : out std_logic;
      total_length_out        : in  integer;
      pcie_bme                : in  std_logic;
      blk_lnk_up              : in  std_logic;
      tag_pending_for_cpl     : in  std_logic;

      -- AXI2PCIE translation vectors
      axibar2pciebar0         : in  std_logic_vector(63 downto 0);
      axibar2pciebar1         : in  std_logic_vector(63 downto 0);
      axibar2pciebar2         : in  std_logic_vector(63 downto 0);
      axibar2pciebar3         : in  std_logic_vector(63 downto 0);
      axibar2pciebar4         : in  std_logic_vector(63 downto 0);
      axibar2pciebar5         : in  std_logic_vector(63 downto 0);
      
      -- AXI Streaming interface
      m_axis_rr_tvalid        : out std_logic;
      m_axis_rr_tready        : in  std_logic;
      m_axis_rr_tdata         : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_rr_tstrb         : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_rr_tlast         : out std_logic;
      config_gen_req          : in  std_logic
   );
end slave_read_req_tlp;

   architecture structure of slave_read_req_tlp is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

--TLP Header Structure

-- Fmt  00      MemWr 3DW (32-bit Address)
--      01      MemWr 4DW (64-bit Address)
-- Type 00000   always for MemRd
-- TC   000     always (default)
-- TD   0       always(no digest field)
-- EP   0       probably won't ever set poison bit
-- Attr 00      always
-- Length       length is inclusive of partial first/last data DWs

-- ReqID        get from PCIe core block IF
-- Tag  x00     not used for MemWr req
-- Last DW BE   generate from ???
-- First DW BE  generate from ???

-- Addr 1 or 2 DW

   type header_array_type is array (0 to 3) of std_logic_vector(31 downto 0);
   signal header_array        : header_array_type;
   signal header_array_reg    : header_array_type;

   type integer_array  is array (0 to 5) of integer range 0 to 1;
   constant C_AXIBAR_AS_ARRAY : integer_array:=(
      C_AXIBAR_AS_0,
      C_AXIBAR_AS_1,
      C_AXIBAR_AS_2,
      C_AXIBAR_AS_3,
      C_AXIBAR_AS_4,
      C_AXIBAR_AS_5);

   type vector_array_type is array (0 to 5) of std_logic_vector(63 downto 0);

   constant C_MASK_ARRAY : vector_array_type := (
                             x"0000_0000_0000_0000" + (C_AXIBAR_0 xor C_AXIBAR_HIGHADDR_0), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_1 xor C_AXIBAR_HIGHADDR_1), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_2 xor C_AXIBAR_HIGHADDR_2), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_3 xor C_AXIBAR_HIGHADDR_3), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_4 xor C_AXIBAR_HIGHADDR_4), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_5 xor C_AXIBAR_HIGHADDR_5));

   constant STR_DATA_SIZE : integer := C_M_AXIS_DATA_WIDTH/32;
   constant FCLIMIT_CPL_V6             : integer := 154*4;
   constant FCLIMIT_CPL_K7             : integer := 154*4;
   constant FCLIMIT_CPL_S6             : integer := 211*4;

   constant FCLIMIT_CPL_FAILSAFE       : integer := 129*4;
   -----------------------------------------------------------------------------
   -- State Machines
   -----------------------------------------------------------------------------

   type rd_req_tlpctlSM_STATES is (IDLE,
                                   SPLIT_REQUEST_1,
                                   SPLIT_REQUEST_2,
                                   SPLIT_REQUEST_3,
                                   BUILD_HEADER,
                                   STR_HEADER_1,
                                   STR_HEADER_2,
                                   STR_HEADER_3,
                                   STR_HEADER_4,
                                   REQ_COMPLETE);
   signal rd_req_tlpctlSM_cs     : rd_req_tlpctlSM_STATES;
   signal rd_req_tlpctlSM_ns     : rd_req_tlpctlSM_STATES;

   signal axibar2pciebar         : vector_array_type;

   signal first_BE               : std_logic_vector(3 downto 0);
   signal first_BE_reg           : std_logic_vector(3 downto 0);
   signal last_BE_reg            : std_logic_vector(3 downto 0);
   signal araddr_2lsbs_reg       : std_logic_vector(1 downto 0);
   signal raddr_reg              : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal rbarhit_reg            : std_logic_vector(C_AXIBAR_NUM-1 downto 0);
   signal length_bytes_reg       : std_logic_vector(12 downto 0);
   signal en_header_array        : std_logic;
   signal enable_addr            : std_logic;
   signal addr_size              : std_logic;
   signal ep                     : std_logic := '0';
   signal address_l              : std_logic_vector(31 downto 0) := x"9ABCDEF0";
   signal address_h              : std_logic_vector(31 downto 0) := x"12345678";
   signal tvalid_int             : std_logic;
   signal tlast_int              : std_logic;
   signal read_req_sent_int      : std_logic;
   signal mrrs_actual            : std_logic_vector(14 downto 0);
   signal first_BE_tmp           : std_logic_vector(3 downto 0);
   signal first_BE_tmp_nxt       : std_logic_vector(3 downto 0);
   signal last_BE_tmp            : std_logic_vector(3 downto 0);
   signal last_BE_tmp_nxt        : std_logic_vector(3 downto 0);
   signal dwlength_tmp           : std_logic_vector(9 downto 0);
   signal dwlength_tmp_nxt       : std_logic_vector(9 downto 0);
   signal dwlength_sent          : std_logic_vector(9 downto 0);
   signal dwlength_sent_nxt      : std_logic_vector(9 downto 0);
   signal address_l_tmp          : std_logic_vector(31 downto 0);
   signal address_l_tmp_nxt      : std_logic_vector(31 downto 0);
   signal num_cmd_splits_nxt     : integer range 0 to 63;
   signal num_cmd_splits         : integer range 0 to 63;
   signal illegal_burst_trns_int : std_logic;
   signal bar_error_trns_int     : std_logic;
   signal tag_count              : integer range 0 to 255;
   signal tag_count_nxt          : integer range 0 to 255;
   signal tag                    : std_logic_vector(7 downto 0) := x"00";
   constant MAX_TAG              : integer range 0 to 255 := 255;
   signal odd_bytes              : integer range 0 to 2;
   signal tlast_d                : std_logic;
   signal fclimit                : integer;
   signal fclimit_block          : std_logic;
   signal s6_limit_adjust        : integer := 0; -- CR # 633509
   signal v6_limit_adjust        : integer := 0; -- CR # 633509
   signal link_down_latch        : std_logic;
   signal first_data_blocked     : std_logic;
   signal v6_limit_adjust_failsafe : integer := 0;

begin

   axibar2pciebar(0)    <= axibar2pciebar0;
   axibar2pciebar(1)    <= axibar2pciebar1;
   axibar2pciebar(2)    <= axibar2pciebar2;
   axibar2pciebar(3)    <= axibar2pciebar3;
   axibar2pciebar(4)    <= axibar2pciebar4;
   axibar2pciebar(5)    <= axibar2pciebar5;
   
   m_axis_rr_tvalid     <= tvalid_int;
   m_axis_rr_tlast      <= tlast_int;
   illegal_burst_trns   <= illegal_burst_trns_int;
   bar_error_trns       <= bar_error_trns_int;

   read_req_sent        <= read_req_sent_int;
   tag_sent             <= tag;

   length_sent          <= dwlength_tmp;
   
   mrrs_actual          <= SHL("000000010000000", maxreadreqsize);
   tag                  <= conv_std_logic_vector(tag_count, 8);

   first_BE               <= x"F" when araddr_2lsbs = "00" and length_bytes > 3 else
                             x"7" when araddr_2lsbs = "00" and length_bytes = 3 else
                             x"3" when araddr_2lsbs = "00" and length_bytes = 2 else
                             x"1" when araddr_2lsbs = "00" and length_bytes = 1 else
                             x"E" when araddr_2lsbs = "01" and length_bytes > 2 else
                             x"6" when araddr_2lsbs = "01" and length_bytes = 2 else
                             x"2" when araddr_2lsbs = "01" and length_bytes = 1 else
                             x"C" when araddr_2lsbs = "10" and length_bytes > 1 else
                             x"4" when araddr_2lsbs = "10" and length_bytes = 1 else
                             x"8";

   address_translation_proccess : process(rbarhit_reg, raddr_reg, axibar2pciebar)
   variable var_addr : std_logic_vector(63 downto 0);
   begin
      var_addr := (others => '0');
      for i in C_AXIBAR_NUM-1 downto 0 loop
         if rbarhit_reg(i) = '1' then
            var_addr := axibar2pciebar(i);
            for j in C_S_AXI_ADDR_WIDTH-1 downto 0 loop
               if(C_MASK_ARRAY(i)(j) = '1') then
                  var_addr(j) := raddr_reg(j);
               end if;
            end loop;
         end if;
         address_l   <= var_addr(31 downto 0);
         address_h   <= var_addr(63 downto 32);
      end loop;
   end process;


   addr_size_proccess : process(rbarhit_reg,axibar2pciebar)
   begin
      addr_size         <= '0';
      for i in C_AXIBAR_NUM-1 downto 0 loop
         if rbarhit_reg(i) = '1' then
            if C_AXIBAR_AS_ARRAY(i) = 1 and axibar2pciebar(i)(63 downto 32) /= x"0000_0000" then
               addr_size         <= '1';
            end if;
         end if;
      end loop;
   end process;


   illegal_burst_trns_proccess : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0' or read_req_sent_int = '1') then
            illegal_burst_trns_int <= '0';
         elsif(illegal_burst = '1') then
            illegal_burst_trns_int <= '1';
         end if;
      end if;
   end process;

   bar_error_trns_proccess : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0' or read_req_sent_int = '1') then
            bar_error_trns_int <= '0';
         elsif(bar_error = '1') then
            bar_error_trns_int <= '1';
         end if;
      end if;
   end process;
   
   odd_bytes_process : process(length_bytes_reg, araddr_2lsbs_reg)
   variable sum : integer;
   begin
      sum := conv_integer(length_bytes_reg(1 downto 0)) + conv_integer(araddr_2lsbs_reg);
      if sum = 0 then
         odd_bytes             <= 0;
      elsif sum < 5 then
         odd_bytes             <= 1;
      else
         odd_bytes             <= 2;
      end if;
   end process;

   s6_limit_adjust <= conv_integer(mrrs_actual(14 downto 2)) when maxreadreqsize(2) = '0' else 256;
   v6_limit_adjust <= conv_integer(mrrs_actual(14 downto 2)) when maxreadreqsize /= "101" else 512;
   
   v6_limit_adjust_failsafe <= 216 when maxreadreqsize = "000" else
                               164 when maxreadreqsize = "001" else
                               conv_integer(mrrs_actual(14 downto 2)) when maxreadreqsize /= "101" else
                               512;
   
   fclimit <= FCLIMIT_CPL_FAILSAFE - v6_limit_adjust_failsafe when C_FAMILY /= "spartan6" and C_EP_LINK_PARTNER_RCB = 0 else
              FCLIMIT_CPL_S6 - s6_limit_adjust when C_FAMILY = "spartan6" else
              FCLIMIT_CPL_V6 - v6_limit_adjust when C_FAMILY = "virtex6" and C_EP_LINK_PARTNER_RCB = 1 else
              FCLIMIT_CPL_K7 - v6_limit_adjust;

   fclimit_block <= '0' when total_length_out < fclimit else '1'; --block requests when fclimit is reached

   link_down_latch_proccess : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            link_down_latch    <= '0';
         elsif link_down_latch = '0' and blk_lnk_up = '0' and
         (tvalid_int = '0' or (tlast_int = '1' and m_axis_rr_tready = '1')) then
            link_down_latch    <= '1';
         elsif(link_down_latch = '1' and blk_lnk_up = '1') then
            link_down_latch    <= '0';
         elsif(first_data_blocked = '1') then
            link_down_latch    <= '1';
         end if;
      end if;
   end process;

   -- This process generates the MemRd TLP(s) that result from one AXI read request
   -- Works with the 'sync' process below 
   rd_req_tlpctlSM_comb : process(rd_req_tlpctlSM_cs, req_active, addr_size, ep, length_bytes_reg, reqID, first_BE_reg,
                                  address_l, address_h, m_axis_rr_tready, mrrs_actual, first_BE_tmp, last_BE_tmp, tag,
                                  dwlength_tmp, address_l_tmp, num_cmd_splits, dwlength_tmp_nxt, last_BE_reg, link_down_latch,
                                  odd_bytes, dwlength_sent, header_array_reg, illegal_burst_trns_int, bar_error_trns_int, fclimit_block,
                                  pcie_bme, blk_lnk_up, tag_pending_for_cpl, config_gen_req)
   begin
      rd_req_tlpctlSM_ns    <= rd_req_tlpctlSM_cs;
      en_header_array       <= '0';
      header_array          <= (others => (others => '0'));
      tlast_int             <= '0';
      m_axis_rr_tdata       <= (others => '0');
      tvalid_int            <= '0';
      m_axis_rr_tstrb       <= (others => '0');
      first_BE_tmp_nxt      <= first_BE_tmp;
      last_BE_tmp_nxt       <= last_BE_tmp;
      dwlength_tmp_nxt      <= dwlength_tmp;
      dwlength_sent_nxt     <= dwlength_sent;
      address_l_tmp_nxt     <= address_l_tmp;
      num_cmd_splits_nxt    <= num_cmd_splits;
      read_req_sent_int     <= '0';
      enable_addr           <= '0';
      first_data_blocked    <= '0';
      case rd_req_tlpctlSM_cs is

         when IDLE =>
            if req_active = '1'  and (pcie_bme = '1' or link_down_latch = '1') then
               enable_addr           <= '1';
               if config_gen_req = '0' then
               rd_req_tlpctlSM_ns    <= SPLIT_REQUEST_1;
	       else
	          rd_req_tlpctlSM_ns    <= IDLE;
	       end if;
            end if;

         when SPLIT_REQUEST_1 =>
            if (length_bytes_reg(12 downto 2) + odd_bytes) <= mrrs_actual(12 downto 2) then
               first_BE_tmp_nxt      <= first_BE_reg;
               dwlength_tmp_nxt      <= length_bytes_reg(11 downto 2) + odd_bytes;
               if dwlength_tmp_nxt = "0000000001" then
                  last_BE_tmp_nxt       <= x"0";
               else
                  last_BE_tmp_nxt       <= last_BE_reg;
               end if;
               address_l_tmp_nxt     <= address_l;
            else--if num_cmd_splits = 0 then
               num_cmd_splits_nxt    <= 1;
               first_BE_tmp_nxt      <= first_BE_reg;
               last_BE_tmp_nxt       <= x"F";
               dwlength_tmp_nxt      <= mrrs_actual(11 downto 2);
               dwlength_sent_nxt     <= mrrs_actual(11 downto 2);
               address_l_tmp_nxt     <= address_l;
            end if;
            rd_req_tlpctlSM_ns    <= BUILD_HEADER;
         when SPLIT_REQUEST_2 =>
            if ((conv_integer(length_bytes_reg(12 downto 2)) + odd_bytes) - dwlength_sent) <= mrrs_actual(12 downto 2)
               then 
               num_cmd_splits_nxt    <= 0;
               dwlength_tmp_nxt      <= (length_bytes_reg(11 downto 2) - dwlength_sent) + odd_bytes;
               rd_req_tlpctlSM_ns    <= SPLIT_REQUEST_3;
            else
               num_cmd_splits_nxt    <= num_cmd_splits + 1;
               first_BE_tmp_nxt      <= x"F";
               last_BE_tmp_nxt       <= x"F";
               dwlength_tmp_nxt      <= mrrs_actual(11 downto 2);
               dwlength_sent_nxt     <= dwlength_sent + mrrs_actual(11 downto 2);
               rd_req_tlpctlSM_ns    <= BUILD_HEADER;
            end if;
            address_l_tmp_nxt     <= address_l_tmp + (dwlength_tmp & "00");

         when SPLIT_REQUEST_3 =>
            if dwlength_tmp = "0000000001" then
               first_BE_tmp_nxt      <= last_BE_reg;
               last_BE_tmp_nxt       <= x"0";
            else
               first_BE_tmp_nxt      <= x"F";
               last_BE_tmp_nxt       <= last_BE_reg;
            end if;
            rd_req_tlpctlSM_ns    <= BUILD_HEADER;

         when BUILD_HEADER =>
            header_array(0)       <= "00" & addr_size & "00" & x"000" & ep & x"0" & dwlength_tmp(9 downto 0);
            header_array(1)       <= reqID & tag & last_BE_tmp & first_BE_tmp;
            if addr_size = '0' then
               header_array(2)       <= address_l_tmp;
               header_array(3)       <= (others => '0');
            else
               header_array(2)       <= address_h;
               header_array(3)       <= address_l_tmp;
            end if;
            if tag_pending_for_cpl = '1' then
              rd_req_tlpctlSM_ns  <= BUILD_HEADER;
            else
              rd_req_tlpctlSM_ns    <= STR_HEADER_1;
            end if;
            en_header_array       <= '1';

         when STR_HEADER_1 =>
            if STR_DATA_SIZE = 1 then    -- 32-bit
               m_axis_rr_tdata    <= header_array_reg(0);
            elsif STR_DATA_SIZE = 2 then -- 64-bit
               m_axis_rr_tdata    <= header_array_reg(1) & header_array_reg(0);
            else--if STR_DATA_SIZE = 4 then -- 128-bit
               tlast_int          <= '1';
               m_axis_rr_tdata    <= header_array_reg(3) & header_array_reg(2) & header_array_reg(1)
                                     & header_array_reg(0);
            end if;
            if illegal_burst_trns_int = '0' and bar_error_trns_int = '0' and fclimit_block = '0' and link_down_latch = '0' and blk_lnk_up = '1' then
               tvalid_int         <= '1';
            end if;
            if STR_DATA_SIZE = 4 then -- 128-bit
               if addr_size = '0' then
                  m_axis_rr_tstrb    <= x"0FFF";
               else
                  m_axis_rr_tstrb    <= (others => '1');
               end if;
            else
               m_axis_rr_tstrb    <= (others => '1');
            end if;
            if (m_axis_rr_tready = '1' and fclimit_block = '0') or illegal_burst_trns_int = '1' or bar_error_trns_int = '1' or link_down_latch = '1' then
               if blk_lnk_up = '0' then
                  first_data_blocked    <= '1';
               end if;
               if STR_DATA_SIZE = 4 then-- 128-bit
                  rd_req_tlpctlSM_ns    <= REQ_COMPLETE;
               else
                  rd_req_tlpctlSM_ns    <= STR_HEADER_2;
               end if;
            end if;

         when STR_HEADER_2 =>
            if STR_DATA_SIZE = 1 then    -- 32-bit
               m_axis_rr_tdata    <= header_array_reg(1);
               -- CR # 646004
            elsif STR_DATA_SIZE = 2 then -- 64-bit
               tlast_int          <= '1';
               m_axis_rr_tdata    <= header_array_reg(3) & header_array_reg(2);
            end if;
            if illegal_burst_trns_int = '0' and bar_error_trns_int = '0' and fclimit_block = '0' and link_down_latch = '0' then
               tvalid_int         <= '1';
            end if;
            if STR_DATA_SIZE = 2 then -- 64-bit
               if addr_size = '0' then 
                  m_axis_rr_tstrb    <= x"0F";
               else
                  m_axis_rr_tstrb    <= (others => '1');
               end if;
            else
               m_axis_rr_tstrb    <= (others => '1');
            end if;
            if (m_axis_rr_tready = '1' and fclimit_block = '0') or illegal_burst_trns_int = '1' or bar_error_trns_int = '1' or link_down_latch = '1' then
               if STR_DATA_SIZE < 2 then
                  rd_req_tlpctlSM_ns    <= STR_HEADER_3;
               else
                  rd_req_tlpctlSM_ns    <= REQ_COMPLETE;
               end if;
            end if;

         when STR_HEADER_3 =>
            m_axis_rr_tdata(31 downto 0)    <= header_array_reg(2);
            if illegal_burst_trns_int = '0' and bar_error_trns_int = '0' and fclimit_block = '0' and link_down_latch = '0' then
               tvalid_int         <= '1';
            end if;
            m_axis_rr_tstrb    <= (others => '1');
            if addr_size = '0' then
               tlast_int          <= '1';
               if (m_axis_rr_tready = '1' and fclimit_block = '0') or illegal_burst_trns_int = '1' or bar_error_trns_int = '1' or link_down_latch = '1' then
                  rd_req_tlpctlSM_ns <= REQ_COMPLETE;
               end if;
            elsif (m_axis_rr_tready = '1' and fclimit_block = '0') or illegal_burst_trns_int = '1' or bar_error_trns_int = '1' or link_down_latch = '1' then
               rd_req_tlpctlSM_ns <= STR_HEADER_4;
            end if;

         when STR_HEADER_4 =>
            m_axis_rr_tdata(31 downto 0)    <= header_array_reg(3);
            if illegal_burst_trns_int = '0' and bar_error_trns_int = '0' and fclimit_block = '0' and link_down_latch = '0' then
               tvalid_int         <= '1';
            end if;
            m_axis_rr_tstrb    <= (others => '1');
            tlast_int          <= '1';
            if (m_axis_rr_tready = '1' and fclimit_block = '0') or illegal_burst_trns_int = '1' or bar_error_trns_int = '1' or link_down_latch = '1' then
               rd_req_tlpctlSM_ns    <= REQ_COMPLETE;
            end if;

         when REQ_COMPLETE =>
            if num_cmd_splits = 0 then
               read_req_sent_int     <= '1';
               rd_req_tlpctlSM_ns    <= IDLE;
            else
               rd_req_tlpctlSM_ns    <= SPLIT_REQUEST_2;
            end if;

      end case;
   end process;

   -- This process generates the MemRd TLP(s) that result from one AXI read request
   -- Works with the 'comb' process above 
   rd_req_tlpctlSM_sync : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            rd_req_tlpctlSM_cs <= IDLE;
            first_BE_tmp       <= (others => '0');
            last_BE_tmp        <= (others => '0');
            dwlength_tmp       <= (others => '0');
            dwlength_sent      <= (others => '0');
            address_l_tmp      <= (others => '0');
            num_cmd_splits     <= 0;
            first_BE_reg       <= (others => '0');
            last_BE_reg        <= (others => '0');
            raddr_reg          <= (others => '0');
            rbarhit_reg        <= (others => '0');
            length_bytes_reg   <= (others => '0');
            header_array_reg   <= (others => (others => '0'));
         else
            rd_req_tlpctlSM_cs <= rd_req_tlpctlSM_ns;
            first_BE_tmp       <= first_BE_tmp_nxt;
            last_BE_tmp        <= last_BE_tmp_nxt;
            dwlength_tmp       <= dwlength_tmp_nxt;
            dwlength_sent      <= dwlength_sent_nxt;
            address_l_tmp      <= address_l_tmp_nxt;
            num_cmd_splits     <= num_cmd_splits_nxt;
            if enable_addr = '1' then
               first_BE_reg       <= first_BE;
               last_BE_reg        <= last_BE;
               raddr_reg          <= raddr;
               rbarhit_reg        <= rbarhit;
               length_bytes_reg   <= length_bytes;
               araddr_2lsbs_reg   <= araddr_2lsbs;
            end if;
            if en_header_array = '1' then
               header_array_reg   <= header_array;
            end if;
         end if;
      end if;
   end process;

-- TAG counter
   tag_counter_comb : process(tag_count, tlast_int, tlast_d)
   begin
      tag_count_nxt         <= tag_count;
      if tlast_int = '0' and tlast_d = '1' then -- neg edge
         if tag_count = MAX_TAG then
            tag_count_nxt         <= 0;
         else
            tag_count_nxt         <= tag_count + 1;
         end if;
      end if;
   end process;

   tag_counter_sync : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            tag_count             <= 0;
            tlast_d               <= '0';
         else
            tag_count             <= tag_count_nxt;
            tlast_d               <= tlast_int;
         end if;
      end if;
   end process;


end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        slave_write_req_tlp.vhd
--
-- Description:     
--                  
-- This VHDL file is an HDL design file for the AXI slave write bridge. 
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              slave_write_req_tlp.vhd
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;


--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------



entity slave_write_req_tlp is
   generic(
      --Family Generics
      C_FAMILY                : string  :="virtex7";

      C_S_AXI_ADDR_WIDTH      : integer := 32;
      C_S_AXI_DATA_WIDTH      : integer := 32;
      C_M_AXIS_DATA_WIDTH     : integer := 32;
      
      C_AXIBAR_NUM            : integer := 6;
      C_AXIBAR_0              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0     : std_logic_vector := x"0000_0000";
      C_AXIBAR_1              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1     : std_logic_vector := x"0000_0000";
      C_AXIBAR_2              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2     : std_logic_vector := x"0000_0000";
      C_AXIBAR_3              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3     : std_logic_vector := x"0000_0000";
      C_AXIBAR_4              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4     : std_logic_vector := x"0000_0000";
      C_AXIBAR_5              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5     : std_logic_vector := x"0000_0000";
      C_AXIBAR_AS_0           : integer := 0;
      C_AXIBAR_AS_1           : integer := 0;
      C_AXIBAR_AS_2           : integer := 0;
      C_AXIBAR_AS_3           : integer := 0;
      C_AXIBAR_AS_4           : integer := 0;
      C_AXIBAR_AS_5           : integer := 0;
      C_AXIBAR_CHK_SLV_ERR    : string  := "FALSE"
   );
   port(

      -- AXI Global
      aclk                    : in  std_logic;
      reset                   : in  std_logic;

      -- internal interface
      maxpayloadsize          : in  std_logic_vector(2 downto 0);
      waddr                   : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      length_bytes            : in  std_logic_vector(12 downto 0);
      wbarhit                 : in  std_logic_vector(C_AXIBAR_NUM-1 downto 0);
      wdata                   : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      first_BE                : in  std_logic_vector(3 downto 0);
      first_BE_valid          : in  std_logic;
      last_BE                 : in  std_logic_vector(3 downto 0);
      last_BE_valid           : in  std_logic;
      first_word_offset       : in  integer;
      wdata_fifo_rd_en        : out std_logic;
      wdata_fifo_empty        : in  std_logic;
      reqID                   : in  std_logic_vector(15 downto 0);
      wdata_str_done          : out std_logic;
      wdata_str_start         : out std_logic;
      illegal_burst_trns      : in  std_logic;
      bar_error_trns          : in  std_logic;
      block_trns_lnkdwn       : in  std_logic;
      blk_lnk_up              : in  std_logic;
      pcie_bme                : in  std_logic;
      tlp_str_start           : out std_logic;

      -- AXI2PCIE translation vectors
      axibar2pciebar0         : in  std_logic_vector(63 downto 0);
      axibar2pciebar1         : in  std_logic_vector(63 downto 0);
      axibar2pciebar2         : in  std_logic_vector(63 downto 0);
      axibar2pciebar3         : in  std_logic_vector(63 downto 0);
      axibar2pciebar4         : in  std_logic_vector(63 downto 0);
      axibar2pciebar5         : in  std_logic_vector(63 downto 0);
      
      -- AXI Streaming interface
      m_axis_rw_tvalid        : out std_logic;
      m_axis_rw_tready        : in  std_logic;
      m_axis_rw_tdata         : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_rw_tstrb         : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_rw_tlast         : out std_logic
      --M_axis_rw_WUSER         : out std_logic_vector()
      
   );
end slave_write_req_tlp;

   architecture structure of slave_write_req_tlp is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

--TLP Header Structure

-- Fmt  10      MemWr 3DW (32-bit Address)
--      11      MemWr 4DW (64-bit Address)
-- Type 00000   always for MemWr
-- TC   000     always (default)
-- TD   0       always(no digest field)
-- EP   0       probably won't ever set poison bit
-- Attr 00      always
-- Length       length is inclusive of partial first/last data DWs

-- ReqID        get from PCIe core block IF
-- Tag  x00     not used for MemWr req
-- Last DW BE   generate from ???
-- First DW BE  generate from ???

-- Addr 1 or 2 DW

   type header_array_type is array (0 to 3) of std_logic_vector(31 downto 0);
   signal header_array        : header_array_type;
   signal header_array_reg    : header_array_type;

   constant ZEROS             : std_logic_vector(127 downto 0) := x"0000_0000_0000_0000_0000_0000_0000_0000";
   constant ONES              : std_logic_vector(15 downto 0) := x"FFFF";
   type integer_array  is array (0 to 5) of integer range 0 to 1;
   constant C_AXIBAR_AS_ARRAY : integer_array:=(
      C_AXIBAR_AS_0,
      C_AXIBAR_AS_1,
      C_AXIBAR_AS_2,
      C_AXIBAR_AS_3,
      C_AXIBAR_AS_4,
      C_AXIBAR_AS_5);

   type vector_array_type is array (0 to 5) of std_logic_vector(63 downto 0);

   constant C_MASK_ARRAY : vector_array_type := (
                             x"0000_0000_0000_0000" + (C_AXIBAR_0 xor C_AXIBAR_HIGHADDR_0), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_1 xor C_AXIBAR_HIGHADDR_1), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_2 xor C_AXIBAR_HIGHADDR_2), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_3 xor C_AXIBAR_HIGHADDR_3), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_4 xor C_AXIBAR_HIGHADDR_4), 
                             x"0000_0000_0000_0000" + (C_AXIBAR_5 xor C_AXIBAR_HIGHADDR_5));

   constant STR_DATA_SIZE : integer := C_M_AXIS_DATA_WIDTH/32;

   -----------------------------------------------------------------------------
   -- State Machines
   -----------------------------------------------------------------------------

   type wr_req_tlpctlSM_STATES is (IDLE,
                                   WAIT_BEs,
                                   WAIT_BME,
                                   SPLIT_REQUEST_1,
                                   SPLIT_REQUEST_2,
                                   SPLIT_REQUEST_3,
                                   LOAD_COUNTER,
                                   BUILD_HEADER,
                                   FIFO_COUNT_ADJ,
                                   STR_HEADER_1,
                                   STR_HEADER_2,
                                   STR_HEADER_3,
                                   STR_HEADER_4,
                                   STR_DATA,
                                   WAIT_BME2);
   signal wr_req_tlpctlSM_cs        : wr_req_tlpctlSM_STATES;
   signal wr_req_tlpctlSM_ns        : wr_req_tlpctlSM_STATES;

   signal axibar2pciebar            : vector_array_type;

   signal first_BE_reg              : std_logic_vector(3 downto 0);
   signal last_BE_reg               : std_logic_vector(3 downto 0);
   signal waddr_reg                 : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal wbarhit_reg               : std_logic_vector(C_AXIBAR_NUM-1 downto 0);
   signal en_header_array           : std_logic;
   signal addr_size                 : std_logic;
   signal ep                        : std_logic := '0';
   signal address_l                 : std_logic_vector(31 downto 0);
   signal address_h                 : std_logic_vector(31 downto 0);
   signal en_data_str               : std_logic;
   signal wdata_fifo_rd_en_int      : std_logic;
   signal wdata_str_done_int        : std_logic;
   signal wdata_str_done_d          : std_logic;
   signal length_bytes_reg          : std_logic_vector(12 downto 0);
   signal fw_offset_reg             : integer;
   signal wr_counter                : integer;
   signal dec_counter               : std_logic;
   signal ld_counter                : std_logic;
   signal wdata_d                   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata_packed              : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal tvalid_int                : std_logic;
   signal tlast_int                 : std_logic;
   signal mps_actual                : std_logic_vector(14 downto 0);
   signal first_BE_tmp              : std_logic_vector(3 downto 0);
   signal first_BE_tmp_nxt          : std_logic_vector(3 downto 0);
   signal last_BE_tmp               : std_logic_vector(3 downto 0);
   signal last_BE_tmp_nxt           : std_logic_vector(3 downto 0);
   signal dwlength_tmp              : std_logic_vector(9 downto 0);
   signal dwlength_tmp_nxt          : std_logic_vector(9 downto 0);
   signal dwlength_sent             : std_logic_vector(9 downto 0);
   signal dwlength_sent_nxt         : std_logic_vector(9 downto 0);
   signal address_l_tmp             : std_logic_vector(31 downto 0);
   signal address_l_tmp_nxt         : std_logic_vector(31 downto 0);
   signal num_cmd_splits_nxt        : integer range 0 to 63;
   signal num_cmd_splits            : integer range 0 to 63;
   signal illegal_burst_latch_int   : std_logic;
   signal bar_error_latch_int       : std_logic;
   signal block_stream_valid        : std_logic;
   signal odd_bytes                 : integer range 0 to 1;
   signal wdata_str_start_int       : std_logic;
   signal block_trns_lnkdwn_latch   : std_logic;
   signal first_data_blocked        : std_logic;
   signal tlp_str_start_int         : std_logic;

-- This function converts a 32-bit little endian format to big endian format
   function little_to_big_endian32(datain : std_logic_vector(31 downto 0))
         return std_logic_vector is
      variable dataout : std_logic_vector(31 downto 0);
   begin
      dataout := datain(7 downto 0) & datain(15 downto 8) & datain(23 downto 16) & datain(31 downto 24);
      return(dataout);
   end function;

begin

   wdata_fifo_rd_en  <= wdata_fifo_rd_en_int;
   m_axis_rw_tvalid  <= tvalid_int;
   m_axis_rw_tlast   <= tlast_int;
   wdata_str_start   <= wdata_str_start_int;
   wdata_str_done    <= wdata_str_done_d;
   tlp_str_start     <= tlp_str_start_int;

   axibar2pciebar(0) <= axibar2pciebar0;
   axibar2pciebar(1) <= axibar2pciebar1;
   axibar2pciebar(2) <= axibar2pciebar2;
   axibar2pciebar(3) <= axibar2pciebar3;
   axibar2pciebar(4) <= axibar2pciebar4;
   axibar2pciebar(5) <= axibar2pciebar5;

   mps_actual <= SHL("000000010000000", maxpayloadsize);

   -- Perform upper bit substitution
   address_translation_proccess : process(wbarhit_reg, waddr_reg, axibar2pciebar)
   variable var_addr : std_logic_vector(63 downto 0);
   begin
      var_addr := (others => '0');
      for i in C_AXIBAR_NUM-1 downto 0 loop
         if wbarhit_reg(i) = '1' then
            var_addr := axibar2pciebar(i);
            for j in C_S_AXI_ADDR_WIDTH-1 downto 0 loop
               if(C_MASK_ARRAY(i)(j) = '1') then
                  var_addr(j) := waddr_reg(j);
               end if;
            end loop;
         end if;
         address_l   <= var_addr(31 downto 0);
         address_h   <= var_addr(63 downto 32);
      end loop;
   end process;


   addr_size_proccess : process(wbarhit_reg,axibar2pciebar)
   begin
      addr_size         <= '0';
      for i in C_AXIBAR_NUM-1 downto 0 loop
         if wbarhit_reg(i) = '1' then
            if C_AXIBAR_AS_ARRAY(i) = 1 and axibar2pciebar(i)(63 downto 32) /= x"0000_0000" then
               addr_size         <= '1';
            end if;
         end if;
      end loop;
   end process;

   illegal_burst_latch_process : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            illegal_burst_latch_int    <= '0';
         elsif(last_BE_valid = '1') then
            illegal_burst_latch_int    <= illegal_burst_trns;
         end if;
      end if;
   end process;

   bar_error_latch_process : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            bar_error_latch_int    <= '0';
         elsif(last_BE_valid = '1') then
            bar_error_latch_int    <= bar_error_trns;
         end if;
      end if;
   end process;

   block_trns_lnkdwn_latch_process : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            block_trns_lnkdwn_latch    <= '0';
         elsif(tlast_int = '1' and m_axis_rw_tready = '1' and block_trns_lnkdwn = '1') -- let current TLP finish, then block
         or (block_trns_lnkdwn = '1' and tvalid_int = '0') -- no TLP, block next
         or (block_trns_lnkdwn = '0' and wdata_str_done_int = '1') -- last TLP blocked, don't block next
         or (block_trns_lnkdwn = '0' and wr_req_tlpctlSM_cs = WAIT_BEs) -- last TLP blocked, don't block next
         then
            block_trns_lnkdwn_latch    <= block_trns_lnkdwn;
         elsif(first_data_blocked = '1') then
            block_trns_lnkdwn_latch    <= '1';
         end if;
      end if;
   end process;

   block_stream_valid <= block_trns_lnkdwn_latch or illegal_burst_latch_int or bar_error_latch_int;

   odd_bytes_process : process(length_bytes_reg)
   begin
      if length_bytes_reg(1 downto 0) /= "00" then
         odd_bytes             <= 1;
      else
         odd_bytes             <= 0;
      end if;
   end process;

   -- This process generates the MemWr TLP(s) that result from one AXI write request, the header is created and streamed
   -- out followed by data from the Write FIFO
   -- Works with the 'sync' and write counter processes below 
   wr_req_tlpctlSM_comb : process(wr_req_tlpctlSM_cs, wbarhit, last_BE_valid, addr_size, ep, length_bytes_reg, reqID,
                                  last_BE_reg, first_BE_reg, address_l, address_h, wdata_fifo_empty, m_axis_rw_tready,
                                  wdata, fw_offset_reg, wr_counter, wdata_packed, mps_actual, first_BE_tmp, last_BE_tmp,
                                  dwlength_tmp, address_l_tmp, num_cmd_splits, dwlength_sent,blk_lnk_up,
                                  header_array_reg, block_stream_valid, odd_bytes, pcie_bme)
   begin
      wr_req_tlpctlSM_ns    <= wr_req_tlpctlSM_cs;
      en_header_array       <= '0';
      header_array          <= (others => (others => '0'));
      wdata_fifo_rd_en_int  <= '0';
      wdata_str_done_int    <= '0';
      wdata_str_start_int   <= '0';
      tlast_int             <= '0';
      en_data_str           <= '0';
      ld_counter            <= '0';
      dec_counter           <= '0';
      m_axis_rw_tdata       <= (others => '0');
      tvalid_int            <= '0';
      m_axis_rw_tstrb       <= (others => '0');
      first_BE_tmp_nxt      <= first_BE_tmp;
      last_BE_tmp_nxt       <= last_BE_tmp;
      dwlength_tmp_nxt      <= dwlength_tmp;
      dwlength_sent_nxt     <= dwlength_sent;
      address_l_tmp_nxt     <= address_l_tmp;
      num_cmd_splits_nxt    <= num_cmd_splits;
      first_data_blocked    <= '0';
      tlp_str_start_int     <= '0';
      case wr_req_tlpctlSM_cs is

         when IDLE =>
            if (C_AXIBAR_CHK_SLV_ERR = "TRUE") then
               wr_req_tlpctlSM_ns <= WAIT_BEs;
            else
               if wbarhit /= ZEROS(C_AXIBAR_NUM-1 downto 0) then-- and (pcie_bme = '1' or block_stream_valid = '1') then
                  wr_req_tlpctlSM_ns <= WAIT_BEs;
               end if;
            end if;

         when WAIT_BEs =>
            if last_BE_valid = '1' then
               wr_req_tlpctlSM_ns    <= WAIT_BME;
            end if;

         when WAIT_BME =>
            -- NAM / JRH fixed typo. Was b 2.
            -- coverage off -item b 1 -allfalse
            if pcie_bme = '1' or block_stream_valid = '1' then
               wr_req_tlpctlSM_ns    <= SPLIT_REQUEST_1;
            end if;

         when SPLIT_REQUEST_1 =>
            if length_bytes_reg <= mps_actual(12 downto 0) then-- less than MPS - no split
               first_BE_tmp_nxt      <= first_BE_reg;
               last_BE_tmp_nxt       <= last_BE_reg;
               dwlength_tmp_nxt      <= length_bytes_reg(11 downto 2) + odd_bytes;
               address_l_tmp_nxt     <= address_l;
            elsif num_cmd_splits = 0 then-- first split
               num_cmd_splits_nxt    <= 1;
               first_BE_tmp_nxt      <= first_BE_reg;
               last_BE_tmp_nxt       <= x"F";
               dwlength_tmp_nxt      <= mps_actual(11 downto 2);
               dwlength_sent_nxt     <= mps_actual(11 downto 2);
               address_l_tmp_nxt     <= address_l;
            end if;
            wr_req_tlpctlSM_ns       <= LOAD_COUNTER;
            tlp_str_start_int        <= '1';

         when SPLIT_REQUEST_2 =>
            if ((conv_integer(length_bytes_reg(11 downto 2)) + odd_bytes) - dwlength_sent) <= mps_actual(11 downto 2)
               then-- last TLP 
               num_cmd_splits_nxt    <= 0;
               dwlength_tmp_nxt      <= (length_bytes_reg(11 downto 2) - dwlength_sent) + odd_bytes;
               wr_req_tlpctlSM_ns    <= SPLIT_REQUEST_3;
            else-- middle TLP
               num_cmd_splits_nxt    <= num_cmd_splits + 1;
               first_BE_tmp_nxt      <= x"F";
               last_BE_tmp_nxt       <= x"F";
               dwlength_tmp_nxt      <= mps_actual(11 downto 2);
               dwlength_sent_nxt     <= dwlength_sent + mps_actual(11 downto 2);
               wr_req_tlpctlSM_ns    <= LOAD_COUNTER;
            end if;
            address_l_tmp_nxt     <= address_l_tmp + (dwlength_tmp & "00");

         when SPLIT_REQUEST_3 =>
            if dwlength_tmp = "0000000001" then
               first_BE_tmp_nxt      <= last_BE_reg;
               last_BE_tmp_nxt       <= x"0";
            else
               first_BE_tmp_nxt      <= x"F";
               last_BE_tmp_nxt       <= last_BE_reg;
            end if;
            wr_req_tlpctlSM_ns    <= LOAD_COUNTER;

         when LOAD_COUNTER =>
            ld_counter            <= '1';
            wr_req_tlpctlSM_ns    <= BUILD_HEADER;

         when BUILD_HEADER =>
            if length_bytes_reg = 0 then
               header_array(0)       <= "01" & addr_size & "00" & x"000" & ep & x"0" & "0000000001";
            else
               header_array(0)       <= "01" & addr_size & "00" & x"000" & ep & x"0" & dwlength_tmp(9 downto 0);
            end if;
            header_array(1)       <= reqID & x"00" & last_BE_tmp & first_BE_tmp;
            if addr_size = '0' then
               header_array(2)       <= address_l_tmp;
               if length_bytes_reg = 0 then -- zero length write TLP
                  header_array(3)    <= (others => '0');
               else
                  header_array(3)    <= little_to_big_endian32(wdata(fw_offset_reg*32+31 downto fw_offset_reg*32));--first_word_offset
                  dec_counter        <= '1';
               end if;
            else
               header_array(2)       <= address_h;
               header_array(3)       <= address_l_tmp;
            end if;
            if (addr_size = '0' or (STR_DATA_SIZE > 1 and fw_offset_reg /= 0)) and length_bytes_reg /= 0 then
               wr_req_tlpctlSM_ns    <= FIFO_COUNT_ADJ;
            else
               wr_req_tlpctlSM_ns    <= STR_HEADER_1;
            end if;
            en_header_array       <= '1';

         when FIFO_COUNT_ADJ =>
            wdata_fifo_rd_en_int  <= '1';
            wr_req_tlpctlSM_ns    <= STR_HEADER_1;

         when STR_HEADER_1 =>
            if num_cmd_splits = 0 then
               wdata_str_start_int   <= '1';
            end if;
            if STR_DATA_SIZE = 1 then    -- 32-bit
               m_axis_rw_tdata       <= header_array_reg(0);
            elsif STR_DATA_SIZE = 2 then -- 64-bit
               m_axis_rw_tdata       <= header_array_reg(1) & header_array_reg(0);
            elsif STR_DATA_SIZE = 4 then -- 128-bit
               m_axis_rw_tdata       <= header_array_reg(3) & header_array_reg(2) & header_array_reg(1)
                                     & header_array_reg(0);
            end if;
            if block_stream_valid = '0' and blk_lnk_up = '1' then
               tvalid_int         <= '1';
            end if;
            m_axis_rw_tstrb    <= (others => '1');
            if STR_DATA_SIZE = 4 then -- 128-bit
               if addr_size = '0' and wr_counter = 0 then
                  tlast_int          <= '1';
                  if m_axis_rw_tready = '1' or block_stream_valid = '1' then
                     if num_cmd_splits = 0 then
                        wr_req_tlpctlSM_ns    <= IDLE;
                        wdata_str_done_int    <= '1';
                        if wdata_fifo_empty = '0' then
                           wdata_fifo_rd_en_int  <= '1';
                        end if;
                     else
                        wr_req_tlpctlSM_ns    <= WAIT_BME2;
                        if(addr_size = '1' and fw_offset_reg = 0 and wdata_fifo_empty = '0') then
                           wdata_fifo_rd_en_int  <= '1';
                        end if;
                     end if;
                  end if;
               elsif m_axis_rw_tready = '1' or block_stream_valid = '1' then
                  wr_req_tlpctlSM_ns    <= STR_DATA;
               end if;
            elsif m_axis_rw_tready = '1' or block_stream_valid = '1' then
               if blk_lnk_up = '0' then
                  first_data_blocked    <= '1';
               end if;
               wr_req_tlpctlSM_ns    <= STR_HEADER_2;
            end if;

         when STR_HEADER_2 =>
            if STR_DATA_SIZE = 1 then    -- 32-bit
               m_axis_rw_tdata    <= header_array_reg(1);
            elsif STR_DATA_SIZE = 2 then -- 64-bit
               m_axis_rw_tdata    <= header_array_reg(3) & header_array_reg(2);
            end if;
            if block_stream_valid = '0' then
               tvalid_int         <= '1';
            end if;
            m_axis_rw_tstrb    <= (others => '1');
            if STR_DATA_SIZE = 2 then
               if addr_size = '0' and wr_counter = 0 then
                  tlast_int          <= '1';
                  if m_axis_rw_tready = '1' or block_stream_valid = '1' then
                     if num_cmd_splits = 0 then
                        wr_req_tlpctlSM_ns    <= IDLE;
                        wdata_str_done_int    <= '1';
                        if wdata_fifo_empty = '0' then
                           wdata_fifo_rd_en_int  <= '1';
                        end if;
                     else
                        wr_req_tlpctlSM_ns    <= WAIT_BME2;
                        if(addr_size = '1' and fw_offset_reg = 0 and wdata_fifo_empty = '0') then
                           wdata_fifo_rd_en_int  <= '1';
                        end if;
                     end if;
                  end if;
               elsif m_axis_rw_tready = '1' or block_stream_valid = '1' then
                  wr_req_tlpctlSM_ns    <= STR_DATA;
               end if;
            elsif m_axis_rw_tready = '1' or block_stream_valid = '1' then
               wr_req_tlpctlSM_ns    <= STR_HEADER_3;
            end if;

         when STR_HEADER_3 =>
            m_axis_rw_tdata(31 downto 0)    <= header_array_reg(2);
            if block_stream_valid = '0' then
               tvalid_int         <= '1';
            end if;
            m_axis_rw_tstrb    <= (others => '1');
            if m_axis_rw_tready = '1' or block_stream_valid = '1' then
               wr_req_tlpctlSM_ns    <= STR_HEADER_4;
            end if;

         when STR_HEADER_4 =>
            m_axis_rw_tdata(31 downto 0)    <= header_array_reg(3);
            if block_stream_valid = '0' then
               tvalid_int         <= '1';
            end if;
            m_axis_rw_tstrb    <= (others => '1');
            if addr_size = '0' and wr_counter = 0 then
               tlast_int          <= '1';
               if m_axis_rw_tready = '1' or block_stream_valid = '1' then
                  if num_cmd_splits = 0 then
                     wr_req_tlpctlSM_ns    <= IDLE;
                     wdata_str_done_int    <= '1';
                     if wdata_fifo_empty = '0' then
                        wdata_fifo_rd_en_int  <= '1';
                     end if;
                  else
                     wr_req_tlpctlSM_ns    <= WAIT_BME2;
                     if(addr_size = '1' and fw_offset_reg = 0 and wdata_fifo_empty = '0') then
                        wdata_fifo_rd_en_int  <= '1';
                     end if;
                  end if;
               end if;
            elsif m_axis_rw_tready = '1' or block_stream_valid = '1' then
               wr_req_tlpctlSM_ns    <= STR_DATA;
            end if;

         when STR_DATA =>
            if block_stream_valid = '0' then
               tvalid_int         <= '1';
            end if;
            if wr_counter < STR_DATA_SIZE and wr_counter /= 0 then
               --m_axis_rw_tdata    <= ZEROS(STR_DATA_SIZE*32-1 downto wr_counter*32)
               --                & wdata_packed(wr_counter*32-1 downto 0);
               --m_axis_rw_tstrb    <= ZEROS(STR_DATA_SIZE*4-1 downto wr_counter*4) & ONES(wr_counter*4-1 downto 0);
               if STR_DATA_SIZE = 2 then -- 64-bit
                  m_axis_rw_tdata    <= ZEROS(63 downto 32)
                                  & wdata_packed(31 downto 0);
                  m_axis_rw_tstrb    <= ZEROS(7 downto 4) & ONES(3 downto 0);
               elsif STR_DATA_SIZE = 4 then -- 128-bit
                  if wr_counter = 3 then
                     m_axis_rw_tdata    <= ZEROS(127 downto 3*32)
                                     & wdata_packed(3*32-1 downto 0);
                     m_axis_rw_tstrb    <= ZEROS(15 downto 3*4) & ONES(3*4-1 downto 0);
                  elsif wr_counter = 2 then
                     m_axis_rw_tdata    <= ZEROS(127 downto 2*32)
                                     & wdata_packed(2*32-1 downto 0);
                     m_axis_rw_tstrb    <= ZEROS(15 downto 2*4) & ONES(2*4-1 downto 0);
                  else
                     m_axis_rw_tdata    <= ZEROS(127 downto 32)
                                     & wdata_packed(31 downto 0);
                     m_axis_rw_tstrb    <= ZEROS(15 downto 4) & ONES(3 downto 0);
                  end if;
               end if;
            else
               if length_bytes_reg = 0 then -- zero length write
                  m_axis_rw_tdata    <= (others => '0');
                  if STR_DATA_SIZE = 1 then -- 32-bit
                     m_axis_rw_tstrb    <= (others => '1');
                  elsif STR_DATA_SIZE = 2 then -- 64-bit
                     m_axis_rw_tstrb    <= ZEROS(7 downto 4) & ONES(3 downto 0);
                  else -- 128-bit
                     m_axis_rw_tstrb    <= ZEROS(15 downto 4) & ONES(3 downto 0);
                  end if;
               else
                  m_axis_rw_tdata    <= wdata_packed;
                  m_axis_rw_tstrb    <= (others => '1');
               end if;
            end if;               
            if wr_counter <= STR_DATA_SIZE then
               tlast_int          <= '1';
               if m_axis_rw_tready = '1' or block_stream_valid = '1' then
                  if num_cmd_splits = 0 then
                     wr_req_tlpctlSM_ns    <= IDLE;
                     wdata_str_done_int    <= '1';
                     if wdata_fifo_empty = '0' then
                        wdata_fifo_rd_en_int  <= '1';
                     end if;
                  else
                     wr_req_tlpctlSM_ns    <= WAIT_BME2;
                     if (STR_DATA_SIZE = 1 or
                     (STR_DATA_SIZE /= 1 and addr_size = '1' and fw_offset_reg = 0))
                     and wdata_fifo_empty = '0' then
                        wdata_fifo_rd_en_int  <= '1';
                     end if;
                  end if;
               end if;
            elsif wdata_fifo_empty = '0' and (m_axis_rw_tready = '1' or block_stream_valid = '1') then
               wdata_fifo_rd_en_int  <= '1';
               en_data_str           <= '1';
            end if;

         when WAIT_BME2 =>
            if pcie_bme = '1' or block_stream_valid = '1' then
               wr_req_tlpctlSM_ns    <= SPLIT_REQUEST_2;
            end if;

      end case;
   end process;

   -- This process generates the MemWr TLP(s) that result from one AXI write request, the header is created and streamed
   -- out followed by data from the Write FIFO
   -- Works with the 'comb' process above and the write counter process below 
   wr_req_tlpctlSM_sync : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            wr_req_tlpctlSM_cs    <= IDLE;
            first_BE_tmp          <= (others => '0');
            last_BE_tmp           <= (others => '0');
            dwlength_tmp          <= (others => '0');
            dwlength_sent         <= (others => '0');
            address_l_tmp         <= (others => '0');
            num_cmd_splits        <= 0;
            wdata_str_done_d      <= '0';
            first_BE_reg          <= (others => '0');
            waddr_reg             <= (others => '0');
            wbarhit_reg           <= (others => '0');
            last_BE_reg           <= (others => '0');
            length_bytes_reg      <= (others => '0');
            fw_offset_reg         <= 0;
            header_array_reg      <= (others => (others => '0'));
         else
            wr_req_tlpctlSM_cs    <= wr_req_tlpctlSM_ns;
            first_BE_tmp          <= first_BE_tmp_nxt;
            last_BE_tmp           <= last_BE_tmp_nxt;
            dwlength_tmp          <= dwlength_tmp_nxt;
            dwlength_sent         <= dwlength_sent_nxt;
            address_l_tmp         <= address_l_tmp_nxt;
            num_cmd_splits        <= num_cmd_splits_nxt;
            wdata_str_done_d      <= wdata_str_done_int;
            if first_BE_valid = '1' then
               first_BE_reg          <= first_BE;
               waddr_reg             <= waddr;
            end if;
            if last_BE_valid = '1' then
               last_BE_reg           <= last_BE;
               length_bytes_reg      <= length_bytes;
               fw_offset_reg         <= first_word_offset;
               wbarhit_reg           <= wbarhit;
            end if;
            if en_header_array = '1' then
               header_array_reg      <= header_array;
            end if;
         end if;
      end if;
   end process;

   wr_counter_proc : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            wr_counter       <= 0;
         else
            if ld_counter = '1' then
               wr_counter       <= conv_integer(dwlength_tmp);
            elsif dec_counter = '1' then
               wr_counter       <= wr_counter-1;
            elsif en_data_str = '1' then
               wr_counter       <= wr_counter-STR_DATA_SIZE;
            end if;
         end if;
      end if;
   end process;

   wdata_delay : process(aclk)
   begin
      if(rising_edge(aclk)) then
         if(reset = '0') then
            wdata_d            <= (others => '0');
         else
            if wdata_fifo_rd_en_int = '1' then
               wdata_d            <= wdata;
            end if;
         end if;
      end if;
   end process;
wdatapacked32: if STR_DATA_SIZE = 1 generate
   data_packer : process(fw_offset_reg, addr_size, wdata, wdata_d)
   begin
         wdata_packed <= little_to_big_endian32(wdata); -- no packing for 32-bit DW
   end process;
end generate wdatapacked32;
wdatapacked64: if STR_DATA_SIZE = 2 generate -- 64-bit
   data_packer : process(fw_offset_reg, addr_size, wdata, wdata_d)
   begin
         if fw_offset_reg = 0 then
            if addr_size = '0' then
               wdata_packed <= little_to_big_endian32(wdata(31 downto 0)) & little_to_big_endian32(wdata_d(63 downto 32)); -- packing for 64-bit DW
            else
               wdata_packed <= little_to_big_endian32(wdata(63 downto 32)) & little_to_big_endian32(wdata(31 downto 0)); -- no packing for 64-bit DW
            end if;
         else -- if fw_offset_reg = 1 then
            if addr_size = '0' then
               wdata_packed <= little_to_big_endian32(wdata(63 downto 32)) & little_to_big_endian32(wdata(31 downto 0)); -- no packing for 64-bit DW
            else
               wdata_packed <= little_to_big_endian32(wdata(31 downto 0)) & little_to_big_endian32(wdata_d(63 downto 32)); -- packing for 64-bit DW
            end if;
         end if;
    end process;
end generate wdatapacked64;
wdatapacked128: if STR_DATA_SIZE = 4 generate -- 128-bit
   data_packer : process(fw_offset_reg, addr_size, wdata, wdata_d)
   begin
         if fw_offset_reg = 0 then
            if addr_size = '0' then
               wdata_packed <=  little_to_big_endian32(wdata(31 downto 0)) & little_to_big_endian32(wdata_d(127 downto 96))
                                & little_to_big_endian32(wdata_d(95 downto 64)) & little_to_big_endian32(wdata_d(63 downto 32)); -- packing for 128-bit DW
            else
               wdata_packed <= little_to_big_endian32(wdata(127 downto 96)) & little_to_big_endian32(wdata(95 downto 64))
                               & little_to_big_endian32(wdata(63 downto 32)) & little_to_big_endian32(wdata(31 downto 0)); -- no packing for 128-bit DW
            end if;
         elsif fw_offset_reg = 1 then
            if addr_size = '0' then
               wdata_packed <= little_to_big_endian32(wdata(63 downto 32)) & little_to_big_endian32(wdata(31 downto 0))
               & little_to_big_endian32(wdata_d(127 downto 96)) & little_to_big_endian32(wdata_d(95 downto 64)); -- packing for 128-bit DW
            else
               wdata_packed <= little_to_big_endian32(wdata(31 downto 0)) & little_to_big_endian32(wdata_d(127 downto 96))
               & little_to_big_endian32(wdata_d(95 downto 64)) & little_to_big_endian32(wdata_d(63 downto 32)); -- packing for 128-bit DW
            end if;
         elsif fw_offset_reg = 2 then
            if addr_size = '0' then
               wdata_packed <= little_to_big_endian32(wdata(95 downto 64)) & little_to_big_endian32(wdata(63 downto 32))
               & little_to_big_endian32(wdata(31 downto 0)) & little_to_big_endian32(wdata_d(127 downto 96)); -- packing for 128-bit DW
            else
               wdata_packed <= little_to_big_endian32(wdata(63 downto 32)) & little_to_big_endian32(wdata(31 downto 0))
               & little_to_big_endian32(wdata_d(127 downto 96)) & little_to_big_endian32(wdata_d(95 downto 64)); -- packing for 128-bit DW
            end if;
         else -- if fw_offset_reg = 3 then
            if addr_size = '0' then
               wdata_packed <= little_to_big_endian32(wdata(127 downto 96)) & little_to_big_endian32(wdata(95 downto 64))
               & little_to_big_endian32(wdata(63 downto 32)) & little_to_big_endian32(wdata(31 downto 0)); -- no packing for 128-bit DW
            else
               wdata_packed <= little_to_big_endian32(wdata(95 downto 64)) & little_to_big_endian32(wdata(63 downto 32))
               & little_to_big_endian32(wdata(31 downto 0)) & little_to_big_endian32(wdata_d(127 downto 96)); -- packing for 128-bit DW
            end if;
         end if;
   end process;
end generate wdatapacked128;
end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_slave_read.vhd
--
-- Description:     
--                  
-- This VHDL file is the HDL design file for the AXI slave write bridge. 
--                   
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_slave_read.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.conv_std_logic_vector;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

entity axi_slave_read is
   generic(
      --Family Generics
      C_FAMILY                      : string  :="virtex7";
      C_S_AXI_ID_WIDTH              : integer := 4;
      C_S_AXI_ADDR_WIDTH            : integer := 32;
      C_S_AXI_DATA_WIDTH            : integer := 32;
      C_COMP_TIMEOUT                : integer := 0; -- 0=50us, 1=50ms
      C_USER_CLK_FREQ               : integer := 1;
      C_USER_CLK2_DIV2              : string  := "FALSE";
      C_S_AXI_SUPPORTS_NARROW_BURST : integer := 1;
      C_AXIREAD_NUM                 : integer := 8;
      C_RD_BUFFER_ADDR_SIZE         : integer := 10;
      C_AXIBAR_NUM                  : integer := 6;
      C_AXIBAR_0                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0           : std_logic_vector := x"0000_0000";
      C_AXIBAR_1                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1           : std_logic_vector := x"0000_0000";
      C_AXIBAR_2                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2           : std_logic_vector := x"0000_0000";
      C_AXIBAR_3                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3           : std_logic_vector := x"0000_0000";
      C_AXIBAR_4                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4           : std_logic_vector := x"0000_0000";
      C_AXIBAR_5                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5           : std_logic_vector := x"0000_0000";
      C_AXIBAR_CHK_SLV_ERR          : string  := "FALSE"
   );
   port(

      -- AXI Global
      s_axi_aclk              : in  std_logic;
      reset                   : in  std_logic;

      -- AXI Slave Read Address Channel
      s_axi_arid              : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_araddr            : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_arregion          : in  std_logic_vector(3 downto 0);
      s_axi_arlen             : in  std_logic_vector(7 downto 0);
      s_axi_arsize            : in  std_logic_vector(2 downto 0);
      s_axi_arburst           : in  std_logic_vector(1 downto 0);
      s_axi_arvalid           : in  std_logic;
      s_axi_arready           : out std_logic;
      pu_axi_arlen            : in  std_logic_vector(7 downto 0);
      pu_axi_arsize           : in  std_logic_vector(2 downto 0);

      -- AXI Slave Read Data Channel
      s_axi_rid               : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_rdata             : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_rresp             : out std_logic_vector(1 downto 0);
      s_axi_rlast             : out std_logic;
      s_axi_rvalid            : out std_logic;
      s_axi_rready            : in  std_logic;

      -- AXIS Read Requester Channel
      m_axis_rr_tid           : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      -- Ordering signals
      slave_read_req_p        : out std_logic;
      slave_rd_req_go         : in  std_logic;
      slave_cmpl_rdy_p        : out std_logic;
      slave_cmpl_go           : in  std_logic;
      slv_write_idle          : in  std_logic;
      master_wr_idle          : in  std_logic;
      -- internal interface
      raddr                   : out std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      length_bytes            : out std_logic_vector(12 downto 0);
      rbarhit                 : out std_logic_vector(C_AXIBAR_NUM-1 downto 0);
      araddr_2lsbs            : out std_logic_vector(1 downto 0);
      last_BE                 : out std_logic_vector(3 downto 0);
      req_active              : out std_logic;
      req_active_ptr          : out integer range 0 to C_AXIREAD_NUM-1;
      read_req_sent           : in  std_logic;
      tag_cpl_status_clr      : in  tag_cpl_status_clr_array;
      rdata_bram_rd_en        : out std_logic;
      rdata_bram_addr         : out std_logic_vector(C_RD_BUFFER_ADDR_SIZE-1 downto 0);
      rdata                   : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      cpl_index               : out integer range 0 to C_AXIREAD_NUM-1;
      rdata_str_done          : out std_logic;
      rdata_str_start         : out std_logic;
      first_word_offset       : out first_word_offset_array;
      illegal_burst           : out std_logic;
      bar_error               : out std_logic;
      cpl_timer_timeout_strb  : out std_logic_vector(C_AXIREAD_NUM-1 downto 0);
      unsupported_req         : in  std_logic;
      completer_abort         : in  std_logic;
      poisoned_req            : in  std_logic_vector(C_AXIREAD_NUM-1 downto 0);
      header_ep               : out std_logic;
      rd_req_index_err        : in  integer range 0 to C_AXIREAD_NUM-1;
      blk_lnk_up              : in  std_logic;
      pcie_bme                : in  std_logic
   );
end axi_slave_read;

architecture structure of axi_slave_read is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

   type addr_array_type is array (natural range <>) of std_logic_vector(31 downto 0);

   constant C_BAR_ADDR_MASK_ARRAY : addr_array_type := (
                             x"0000_0000" + C_AXIBAR_0 xnor C_AXIBAR_HIGHADDR_0, 
                             x"0000_0000" + C_AXIBAR_1 xnor C_AXIBAR_HIGHADDR_1, 
                             x"0000_0000" + C_AXIBAR_2 xnor C_AXIBAR_HIGHADDR_2, 
                             x"0000_0000" + C_AXIBAR_3 xnor C_AXIBAR_HIGHADDR_3, 
                             x"0000_0000" + C_AXIBAR_4 xnor C_AXIBAR_HIGHADDR_4, 
                             x"0000_0000" + C_AXIBAR_5 xnor C_AXIBAR_HIGHADDR_5);

   constant C_BAR_HIGHADDR_ARRAY : addr_array_type := (C_AXIBAR_HIGHADDR_0, 
                                                       C_AXIBAR_HIGHADDR_1, 
                                                       C_AXIBAR_HIGHADDR_2, 
                                                       C_AXIBAR_HIGHADDR_3, 
                                                       C_AXIBAR_HIGHADDR_4, 
                                                       C_AXIBAR_HIGHADDR_5);

   constant C_BAR_ARRAY : addr_array_type := (C_AXIBAR_0, 
                                              C_AXIBAR_1, 
                                              C_AXIBAR_2, 
                                              C_AXIBAR_3, 
                                              C_AXIBAR_4, 
                                              C_AXIBAR_5);

   constant DATA_SIZE                  : integer := C_S_AXI_DATA_WIDTH/32;
   constant HISTORY_SIZE               : integer := C_AXIREAD_NUM;

   constant ONES                       : std_logic_vector(0 to DATA_SIZE*8-1) := (others => '1');
   constant ZEROES                     : std_logic_vector(0 to DATA_SIZE*8-1) := (others => '0');
   type arid_array is array (0 to C_AXIREAD_NUM-1) of std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
   signal arid_reg                     : arid_array := (others => (others => '0'));  -- CR # 649227
   signal araddr_reg                   : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal arregion_reg                 : std_logic_vector(3 downto 0);
   type arlen_array is array (0 to C_AXIREAD_NUM-1) of std_logic_vector(7 downto 0);
   signal arlen_reg                    : arlen_array;
   --signal arsize_reg                   : std_logic_vector(2 downto 0);
   signal arburst_reg                  : std_logic_vector(1 downto 0);
   signal rd_req_ptr                   : integer range 0 to C_AXIREAD_NUM-1 := 0;
   signal rd_req_ptr_nxt               : integer range 0 to C_AXIREAD_NUM-1 := 0;
   type arid_history_array is array (0 to HISTORY_SIZE-1) of std_logic_vector(C_S_AXI_ID_WIDTH downto 0);
   signal arid_history                 : arid_history_array;
   signal arid_history_nxt             : arid_history_array;
   type rd_req_ptr_array is array (0 to HISTORY_SIZE-1) of integer range 0 to C_AXIREAD_NUM-1;
   signal rd_req_ptr_history           : rd_req_ptr_array;
   signal rd_req_ptr_history_nxt       : rd_req_ptr_array;
   constant ZEROS                      : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  -- constant ZEROS                      : std_logic_vector(12 downto 0) := "0000000000000";
   signal barhit                       : std_logic_vector(C_AXIBAR_NUM-1 downto 0);
   signal arready_int                  : std_logic;
   signal s_axi_rlast_int              : std_logic := '0';  -- CR # 649227
   signal s_axi_rdata_int              : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0) := (others => '0');  -- CR # 649227
   signal s_axi_rresp_int              : std_logic_vector(1 downto 0) := (others => '0');  -- CR # 649227
   signal rvalid_int                   : std_logic := '0';
   signal illegal_burst_int            : std_logic;
   signal bar_error_int                : std_logic;
   signal read_req_error               : std_logic;
   signal en_barhit                    : std_logic;
   signal rlast_int                    : std_logic := '0';
   signal en_rresp                     : std_logic := '0';
   signal size                         : integer range 1 to 16;
   signal length_bytes_int             : std_logic_vector(12 downto 0);
   signal first_word_offset_int        : first_word_offset_array;
   signal first_word_offset_calc       : integer range 0 to 3;
   signal rdata_bram_rd_en_int         : std_logic;
   signal rd_counter                   : integer range 0 to 511;
   signal rdata_str_done_int           : std_logic;
   signal rd_req_index                 : integer range 0 to C_AXIREAD_NUM-1 := 0;
   signal cpl_index_int                : integer range 0 to C_AXIREAD_NUM-1;
   signal cpl_index_nxt                : integer range 0 to C_AXIREAD_NUM-1;
   signal open_slot                    : std_logic;
   signal slot_cleared                 : std_logic;
   signal slot_cleared_d               : std_logic;
   signal slot_request                 : std_logic;
   signal pending_rd_reqs              : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal pending_rd_reqs_nxt          : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal pending_rd_reqs_d            : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal pu_arlen_reg                 : std_logic_vector(7 downto 0);
   signal pu_arsize_reg                : std_logic_vector(2 downto 0);
   signal pu_length_bytes              : std_logic_vector(12 downto 0);
   signal arid_match_index             : integer range 0 to HISTORY_SIZE-1;
   signal arid_match_index_nxt         : integer range 0 to HISTORY_SIZE-1;
   signal dependency_ptr               : integer range 0 to C_AXIREAD_NUM-1;
   type arid_dependency_array is array (0 to C_AXIREAD_NUM-1) of integer range 0 to C_AXIREAD_NUM;
   signal arid_dependency              : arid_dependency_array;
   signal arid_dependency_nxt          : arid_dependency_array;
   type arid_rresp_array is array (0 to C_AXIREAD_NUM-1) of std_logic_vector(1 downto 0);
   signal arid_rresp                   : arid_rresp_array := (others => (others => '0'));  -- CR # 649227
   signal new_dependency_entry         : std_logic;
   signal clr_dependency_entry         : std_logic;
   signal new_dependency_hs            : std_logic;
   signal dependency_cleared           : std_logic;
   signal no_pending_reqs              : std_logic;
   signal clr_pending_rd_reqs_entry    : std_logic;
   signal rdata_mask                   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal cpl_timer_start_count        : integer;
   signal tag_cpl_status_clr_d         : tag_cpl_status_clr_array;
   type cpl_timer_count_array is array (0 to C_AXIREAD_NUM-1,0 to C_S_AXI_DATA_WIDTH/4-1) of integer range 0 to (2**14 + ((2**24)-(2**14))*C_COMP_TIMEOUT) - 1;
   signal cpl_timer_count              : cpl_timer_count_array;
   signal cpl_timer_count_nxt          : cpl_timer_count_array;
   signal cpl_timer_timeout            : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal cpl_timer_timeout_int        : tag_cpl_status_clr_array;
   signal cpl_timer_timeout_d          : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal cpl_timer_timeout_strb_int   : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal blk_lnk_up_d                 : std_logic;
   signal cpl_req_index                : integer range 0 to C_AXIREAD_NUM;
   signal cpl_permit                   : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal req_active_int               : std_logic;
   signal ld_rd_counter                : std_logic;
   signal slv_rd_req_p_sent            : std_logic;
   signal slave_cmpl_go_pend           : std_logic;
   signal cmpl_rdy_pend                : std_logic_vector(C_AXIREAD_NUM-1 downto 0);

   -----------------------------------------------------------------------------
   -- State Machines
   -----------------------------------------------------------------------------

   type read_reqSM_STATES is (IDLE,
                              CHECK,
                              SEND_REQ,
                              WAIT_FOR_OPEN_SLOT);
   signal read_reqSM_cs : read_reqSM_STATES;
   signal read_reqSM_ns : read_reqSM_STATES;

   type read_dataSM_STATES is (IDLE,
                               WAIT_FOR_CPL,
                               LOAD_READ_COUNTER,
                               FIRST_BRAM_READ,
                               STR_DATA,
                               STR_DONE,
                               WAIT_SLOT_CLR);
   signal read_dataSM_cs : read_dataSM_STATES;
   signal read_dataSM_ns : read_dataSM_STATES;
   signal read_dataSM_cs_d : read_dataSM_STATES;
   
   type arid_dependencySM_STATES is (IDLE,
                                     FIND_HISTORY_MATCH,
                                     SET_DEPENDENCY,
                                     CLEAR_DEPENDENCY);
   signal arid_dependencySM_cs : arid_dependencySM_STATES;
   signal arid_dependencySM_ns : arid_dependencySM_STATES;
   
begin

   s_axi_rlast            <= s_axi_rlast_int;  -- CR # 649227
   s_axi_rdata            <= s_axi_rdata_int;   -- CR # 649227
   s_axi_rresp            <= s_axi_rresp_int;  -- CR # 649227
   s_axi_arready          <= arready_int;
   s_axi_rvalid           <= rvalid_int;
   illegal_burst          <= illegal_burst_int;
   bar_error              <= bar_error_int;
   s_axi_rid              <= arid_reg(cpl_index_int);
   m_axis_rr_tid          <= arid_reg(rd_req_ptr);
   cpl_timer_timeout_strb <= cpl_timer_timeout_strb_int;

   -- CR # 649227
   s_axi_rresp_int        <= arid_rresp(cpl_index_int) when en_rresp = '1' and (blk_lnk_up = '1' or
                                                           (blk_lnk_up = '0'and read_dataSM_cs_d = STR_DATA))
                             else
                             "10"  when en_rresp = '1' and blk_lnk_up = '0' and read_dataSM_cs_d = FIRST_BRAM_READ -- SLVERR
                             else (others => '0');

   req_active_ptr         <= rd_req_ptr;
   req_active             <= req_active_int;
   rdata_str_done         <= rdata_str_done_int;
   cpl_index              <= cpl_index_int;
   araddr_2lsbs           <= araddr_reg(1 downto 0);
   first_word_offset      <= first_word_offset_int;

   -- Generate the read buffer address for getting read return data to the AXI4
   rdata_bram_addr        <= conv_std_logic_vector(cpl_index_int, log2(C_AXIREAD_NUM))
                             & conv_std_logic_vector(conv_integer(arlen_reg(cpl_index_int)) - rd_counter + 1, 8);
   rdata_bram_rd_en       <= rdata_bram_rd_en_int;


   length_bytes           <= pu_length_bytes;

   pu_length_bytes        <= ("00000" & pu_arlen_reg) + 1 when pu_arsize_reg = "000"
                             else
                             --SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto conv_integer(pu_arsize_reg)) & araddr_reg(conv_integer(pu_arsize_reg)
                             -- - 1 downto 0));
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 1) & araddr_reg(0 downto 0)) when pu_arsize_reg = "001" else
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 2) & araddr_reg(1 downto 0)) when pu_arsize_reg = "010" else
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 3) & araddr_reg(2 downto 0)) when pu_arsize_reg = "011" else
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 4) & araddr_reg(3 downto 0)) when pu_arsize_reg = "100" else
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 5) & araddr_reg(4 downto 0)) when pu_arsize_reg = "101" else
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 6) & araddr_reg(5 downto 0)) when pu_arsize_reg = "110" else
                             SHL(("00000" & pu_arlen_reg) + 1, pu_arsize_reg) - (ZEROS(12 downto 7) & araddr_reg(6 downto 0));

   last_BE                <= x"1" when (conv_integer(araddr_reg(1 downto 0)) + conv_integer(pu_length_bytes(1 downto 0)))
                                       mod 4 = 1 else
                             x"3" when (conv_integer(araddr_reg(1 downto 0)) + conv_integer(pu_length_bytes(1 downto 0)))
                                       mod 4 = 2 else
                             x"7" when (conv_integer(araddr_reg(1 downto 0)) + conv_integer(pu_length_bytes(1 downto 0)))
                                       mod 4 = 3 else
                             x"F";

   first_word_offset_calc <= 0 when DATA_SIZE = 1 or (DATA_SIZE = 2 and s_axi_araddr(2) = '0') or
                                    (DATA_SIZE = 4 and s_axi_araddr(3 downto 2) = "00") else
                             1 when (DATA_SIZE = 2 and s_axi_araddr(2) = '1') or
                                    (DATA_SIZE = 4 and s_axi_araddr(3 downto 2) = "01") else
                             2 when (DATA_SIZE = 4 and s_axi_araddr(3 downto 2) = "10") else
                             3;

   raddr                  <= araddr_reg(C_S_AXI_ADDR_WIDTH-1 downto 2) & "00"
                                when first_word_offset_int(rd_req_ptr) = 0
                             else araddr_reg(C_S_AXI_ADDR_WIDTH-1 downto 3) & "100"
                                when first_word_offset_int(rd_req_ptr) = 1
                             else araddr_reg(C_S_AXI_ADDR_WIDTH-1 downto 4) & "1000"
                                when first_word_offset_int(rd_req_ptr) = 2
                             else araddr_reg(C_S_AXI_ADDR_WIDTH-1 downto 4) & "1100";

   gen_rdata_mask_32 : if C_S_AXI_DATA_WIDTH = 32 generate
      rdata_mask             <= (others => '1') after 100 ps;
   end generate;

   gen_rdata_mask_64 : if C_S_AXI_DATA_WIDTH = 64 generate
      rdata_mask             <= x"FFFF_FFFF_0000_0000"  after 100 ps when rd_counter = conv_integer(arlen_reg(cpl_index_int)) and
                                first_word_offset_int(cpl_index_int) = 1
                             else
                             (others => '1') after 100 ps;
   end generate;

   gen_rdata_mask_128 : if C_S_AXI_DATA_WIDTH = 128 generate
      rdata_mask             <= x"FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_0000_0000"  after 100 ps when rd_counter = conv_integer(arlen_reg(cpl_index_int))
                                and first_word_offset_int(cpl_index_int) = 1
                             else
                             x"FFFF_FFFF_FFFF_FFFF_0000_0000_0000_0000"  after 100 ps when rd_counter = conv_integer(arlen_reg(cpl_index_int))
                                and first_word_offset_int(cpl_index_int) = 2
                             else
                             x"FFFF_FFFF_0000_0000_0000_0000_0000_0000"  after 100 ps when rd_counter = conv_integer(arlen_reg(cpl_index_int))
                                and first_word_offset_int(cpl_index_int) = 3
                             else
                             (others => '1') after 100 ps;
   end generate;

   slv_rd_req_p_sent_proccess :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0' or req_active_int = '1') then
            slv_rd_req_p_sent            <= '0';
         elsif s_axi_arvalid = '1' and arready_int = '1' and slv_write_idle = '0' then
            slv_rd_req_p_sent            <= '1';
         end if;
      end if;
   end process;

   gen_cpl_timer_timeout : for j in 0 to C_AXIREAD_NUM-1 generate
      cpl_timer_timeout(j) <= '0' when cpl_timer_timeout_int(j)(0 to DATA_SIZE*8-1) = ZEROES else '1';
   end generate gen_cpl_timer_timeout;

   -- Get read address phase info from AXI for up to 8 "slots" when available
   -- Works with the 'sync' process below 
   read_reqSM_comb :process(read_reqSM_cs, s_axi_arvalid, barhit, read_req_sent, open_slot, rd_req_ptr, blk_lnk_up,
                            arburst_reg, arid_rresp, slave_rd_req_go, slv_rd_req_p_sent, pcie_bme)
   begin
      read_reqSM_ns          <= read_reqSM_cs;
      arready_int            <= '0';
      req_active_int         <= '0';
      illegal_burst_int      <= '0';
      bar_error_int          <= '0';
      en_barhit              <= '0';
      read_req_error         <= '0';
      slot_request           <= '0';
      case read_reqSM_cs is

         when IDLE =>
            if blk_lnk_up = '1' and pcie_bme = '1' then -- only assert awready if link is up
               arready_int         <= '1';
            end if;
            if s_axi_arvalid = '1' and blk_lnk_up = '1' and pcie_bme = '1' then
               -- aquire read req qualifiers
               read_reqSM_ns       <= CHECK;
            end if;

         when CHECK =>
            -- check qualifiers
            en_barhit           <= '1';
            -- coverage off
            -- never hit, remove in 13.3
            if barhit = ZEROS(C_AXIBAR_NUM - 1 downto 0) then
               if (C_AXIBAR_CHK_SLV_ERR = "TRUE") then
                  bar_error_int       <= '1';
                  read_reqSM_ns       <= SEND_REQ;
               else
                  bar_error_int       <= '0';
                  read_reqSM_ns       <= IDLE;
               end if;
            -- coverage on
            elsif slave_rd_req_go = '1' or slv_rd_req_p_sent = '0' or blk_lnk_up = '0' then
               read_reqSM_ns       <= SEND_REQ;
            end if;
            if (arburst_reg /= "01") then
               illegal_burst_int   <= '1';
               read_reqSM_ns       <= SEND_REQ;
            end if;

         when SEND_REQ =>
            req_active_int      <= '1';
            if read_req_sent = '1' then
               read_reqSM_ns       <= WAIT_FOR_OPEN_SLOT;
            end if;

         when WAIT_FOR_OPEN_SLOT =>
            slot_request        <= '1';
            if open_slot = '1' then
               read_reqSM_ns       <= IDLE;
            end if;

      end case;
   end process;

   -- Get read address phase info from AXI for up to 8 "slots" when available
   -- Works with the 'comb' process above 
   read_reqSM_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            read_reqSM_cs                <= IDLE;
            arid_reg                     <= (others => (others => '0'));
            araddr_reg                   <= (others => '0');
            arregion_reg                 <= (others => '0');
            arlen_reg                    <= (others => (others => '0'));
            arburst_reg                  <= (others => '0');
            pu_arlen_reg                 <= (others => '0');
            pu_arsize_reg                <= (others => '0');
            rbarhit                      <= (others => '0');
            first_word_offset_int        <= (others => 0);
            slave_read_req_p             <= '0';
         else
            read_reqSM_cs <= read_reqSM_ns;
            slave_read_req_p             <= '0';
            if s_axi_arvalid = '1' and arready_int = '1' then
               arid_reg(rd_req_ptr)         <= s_axi_arid;
               araddr_reg                   <= s_axi_araddr;
               arregion_reg                 <= s_axi_arregion;
               arlen_reg(rd_req_ptr)        <= s_axi_arlen;
               arburst_reg                  <= s_axi_arburst;
               pu_arlen_reg                 <= pu_axi_arlen; --pu means pre-upsizer
               pu_arsize_reg                <= pu_axi_arsize;
               first_word_offset_int(rd_req_ptr)   <= first_word_offset_calc;
               slave_read_req_p             <= not(slv_write_idle);
            end if;
            if en_barhit = '1' then
               rbarhit             <= barhit;
            end if;
         end if;
      end if;
   end process;

   BAR_decoder :process(araddr_reg)

--   Remove the use of ARRegion
--   BAR_decoder :process(arregion_reg)
--   variable region    : integer;
--
--   begin
--      region                 := conv_integer(arregion_reg);
--      barhit                 <= (others => '0');
--      -- Nam - always true if statement below
--      -- NAM / JRH fixed typo. Was b 2.
--      -- coverage off -item b 1 -allfalse
--      if region < C_AXIBAR_NUM then
--         barhit(region)         <= '1';
--      end if;
   variable address : integer;
   begin
--     address := conv_integer(araddr_reg);
     barhit <= (others => '0');

     -- Nam - always true if statement below
     -- NAM /JRH fixed typo. Was b 2.
     -- coverage off -item b 1 -allfalse
     for i in 0 to (C_AXIBAR_NUM-1) loop
       if((araddr_reg <= C_BAR_HIGHADDR_ARRAY(i)) and (araddr_reg >= C_BAR_ARRAY(i))) then
         barhit(i) <= '1';
       end if;
     end loop;       
   end process;

   -- This process maintains the pending read status vector of 8 'slots' for AXI read requests
   -- Works with the 'sync' process below 
   pend_rdreq_status_comb :process(read_req_sent, illegal_burst_int, bar_error_int, slot_request, clr_pending_rd_reqs_entry, arid_reg,
                                   pending_rd_reqs, cpl_index_int, rd_req_ptr, arid_history, rd_req_ptr_history)
   variable first_zero  : boolean;
   variable first_match : boolean;
   variable index_save  : integer range 0 to HISTORY_SIZE;
   variable clear_mask8 : unsigned(0 to HISTORY_SIZE-1);-- := x"FE";
   variable clear_mask4 : unsigned(0 to 3) := x"E";
   begin
      if HISTORY_SIZE = 8 then
         clear_mask8 := x"FE";
      else
         clear_mask8 := x"E";
      end if;
      rd_req_ptr_nxt         <= rd_req_ptr;
      pending_rd_reqs_nxt    <= pending_rd_reqs;
      open_slot              <= '0';
      slot_cleared           <= '0';
      arid_history_nxt       <= arid_history;
      rd_req_ptr_history_nxt <= rd_req_ptr_history;
      if read_req_sent = '1' then
         if HISTORY_SIZE = 8 then
            pending_rd_reqs_nxt    <= pending_rd_reqs or SHL(x"01", conv_std_logic_vector(rd_req_ptr, 3));
         else
            pending_rd_reqs_nxt    <= pending_rd_reqs or SHL(x"1", conv_std_logic_vector(rd_req_ptr, 2));
         end if;
         arid_history_nxt       <= ('1' & arid_reg(rd_req_ptr)) & arid_history(0 to HISTORY_SIZE-2);
         rd_req_ptr_history_nxt <= rd_req_ptr & rd_req_ptr_history(0 to HISTORY_SIZE-2);
      elsif clr_pending_rd_reqs_entry = '1' then -- clear pending read request
         pending_rd_reqs_nxt    <= pending_rd_reqs and STD_LOGIC_VECTOR(rotate_left(clear_mask8, cpl_index_int));
         slot_cleared           <= '1';
         first_match            := FALSE;
         for i in 0 to HISTORY_SIZE-1 loop -- find the most recent pending read request of current arid
            if rd_req_ptr_history(i) = cpl_index_int and--arid_history(i)(C_S_AXI_ID_WIDTH) = '1' and
            first_match = FALSE then
               first_match            := TRUE;
               arid_history_nxt(i to HISTORY_SIZE-1) <= arid_history(i+1 to HISTORY_SIZE-1)
                                                        & ZEROS(C_S_AXI_ID_WIDTH downto 0);
               rd_req_ptr_history_nxt(i to HISTORY_SIZE-2) <= rd_req_ptr_history(i+1 to HISTORY_SIZE-1);
            end if;
         end loop;
      elsif slot_request = '1' then
         first_zero             := FALSE;
         index_save             := HISTORY_SIZE;
         for i in 0 to C_AXIREAD_NUM-1 loop -- find lowest open read request slot
            if pending_rd_reqs(i) = '0' and first_zero = FALSE then
               first_zero             := TRUE;
               index_save             := i;
            end if;
         end loop;
         if index_save /= HISTORY_SIZE then -- set pending read request
            open_slot              <= '1';
            rd_req_ptr_nxt         <= index_save;
         end if;
      end if;
   end process;

   -- This process maintains the pending read status vector of 8 'slots' for AXI read requests
   -- Works with the 'comb' process above 
   pend_rdreq_status_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            pending_rd_reqs        <= (others => '0');
            pending_rd_reqs_d      <= (others => '0');
            rd_req_ptr             <= 0;
            arid_history           <= (others => (others => '0'));
            rd_req_ptr_history     <= (others => 0);
            clr_pending_rd_reqs_entry          <= '0';
            slot_cleared_d         <= '0';
         else
            pending_rd_reqs        <= pending_rd_reqs_nxt;
            pending_rd_reqs_d      <= pending_rd_reqs;
            rd_req_ptr             <= rd_req_ptr_nxt;
            arid_history           <= arid_history_nxt;
            rd_req_ptr_history     <= rd_req_ptr_history_nxt;
            slot_cleared_d         <= slot_cleared;
            if rdata_str_done_int = '1' then
               clr_pending_rd_reqs_entry          <= '1';
            elsif slot_cleared_d = '1' then
               clr_pending_rd_reqs_entry          <= '0';
            end if;
         end if;
      end if;
   end process;


   -- This process maintains the 'slot' buffer data dependencies that are an array of integer values that are assigned
   -- values N as follows:
   -- N = 8 for no dependency, N = 0 - 7 indicates dependency on 'slot' buffer N
   -- Works with the 'sync' process below 
   arid_dependencySM_comb :process(arid_dependencySM_cs, new_dependency_entry, arid_history, rd_req_ptr_history, arid_reg,
                                   arid_match_index, arid_dependency, dependency_ptr, pending_rd_reqs, no_pending_reqs,
                                   clr_dependency_entry, cpl_index_int, clr_pending_rd_reqs_entry)
   variable first_match  : boolean;
   begin
      arid_dependencySM_ns                  <= arid_dependencySM_cs;
      arid_match_index_nxt                  <= arid_match_index;
      arid_dependency_nxt                   <= arid_dependency;  
      new_dependency_hs                     <= '0';
      dependency_cleared                    <= '0';
      case arid_dependencySM_cs is
         when IDLE =>
            if clr_dependency_entry = '1' then
               arid_dependencySM_ns   <= CLEAR_DEPENDENCY;
            elsif new_dependency_entry = '1' and clr_pending_rd_reqs_entry = '0' then
               arid_dependencySM_ns   <= FIND_HISTORY_MATCH;
            end if;

         when FIND_HISTORY_MATCH =>
            if clr_pending_rd_reqs_entry = '0' then
               if C_S_AXI_SUPPORTS_NARROW_BURST = 0 then -- use arid matching for multi thread
                  first_match            := FALSE;
                  for i in 1 to HISTORY_SIZE-1 loop -- find the most recent pending read request of current arid
                     if arid_history(i) = ('1' & arid_reg(dependency_ptr)) and pending_rd_reqs(rd_req_ptr_history(i)) = '1'
                     and first_match = FALSE then
                        first_match            := TRUE;
                        arid_match_index_nxt   <= i;
                     end if;
                  end loop;
               elsif no_pending_reqs = '0' then -- don't use arid matching for multi thread
                  if arid_history(1)(C_S_AXI_ID_WIDTH) = '1' then
                     first_match            := TRUE;
                     arid_match_index_nxt   <= 1;
                  else
                     first_match            := FALSE;
                  end if;
               else
                  first_match            := FALSE;
               end if;
               if first_match = TRUE then
                  arid_dependencySM_ns                  <= SET_DEPENDENCY;
               else
                  arid_dependencySM_ns                  <= IDLE;
                  new_dependency_hs                     <= '1';
               end if;
            end if;

         when SET_DEPENDENCY =>
            if pending_rd_reqs(rd_req_ptr_history(arid_match_index)) = '1' then -- match is still pending
               arid_dependency_nxt(dependency_ptr)   <= rd_req_ptr_history(arid_match_index);
            else
               arid_dependency_nxt(dependency_ptr)   <= HISTORY_SIZE;
            end if;
            arid_dependencySM_ns                  <= IDLE;
            new_dependency_hs                     <= '1';

         when CLEAR_DEPENDENCY =>
            first_match                           := FALSE;
            for i in 0 to C_AXIREAD_NUM-1 loop --find and clear dependency on this completion
               if arid_dependency(i) = cpl_index_int and first_match = FALSE then
                  first_match                           := TRUE;
                  arid_dependency_nxt(i)                <= HISTORY_SIZE;
               end if;
            end loop;
            dependency_cleared                    <= '1';
            arid_dependencySM_ns                  <= IDLE;

      end case;
   end process;

   -- This process maintains the 'slot' buffer data dependencies that are an array of integer values that are assigned
   -- values N as follows:
   -- N = 8 for no dependency, N = 0 - 7 indicates dependency on 'slot' buffer N
   -- Works with the 'comb' process above 
   arid_dependencySM_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            arid_dependencySM_cs               <= IDLE;
            arid_dependency                    <= (others => HISTORY_SIZE);
            arid_match_index                   <= 0;
            dependency_ptr                     <= 0;
            new_dependency_entry               <= '0';
            clr_dependency_entry               <= '0';
            no_pending_reqs                    <= '0';
         else
            arid_dependencySM_cs               <= arid_dependencySM_ns;
            arid_dependency                    <= arid_dependency_nxt;
            arid_match_index                   <= arid_match_index_nxt;
            if read_req_sent = '1' then
               dependency_ptr                     <= rd_req_ptr;
               new_dependency_entry               <= '1';
               if HISTORY_SIZE = 8 then
                  if pending_rd_reqs = x"00" then
                     no_pending_reqs                    <= '1';
                  end if;
               else
                  if pending_rd_reqs = x"0" then
                     no_pending_reqs                    <= '1';
                  end if;
               end if;
            elsif new_dependency_hs = '1' then
               new_dependency_entry               <= '0';
               no_pending_reqs                    <= '0';
            end if;
            if rdata_str_done_int = '1' then
               clr_dependency_entry               <= '1';
            elsif dependency_cleared = '1' then
               clr_dependency_entry               <= '0';
            end if;
         end if;
      end if;
   end process;

   -- This process maintains rresp for each 'slot' read request
   -- After each 'slot' buffer is read and data returned to the AXI read channel, the 'slot' rresp value is cleared
   -- Different error conditions will set the 'slot' rresp value to SLVERR
   rresp_gen :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            arid_rresp         <= (others => (others => '0')); -- OKAY is default
            blk_lnk_up_d       <= '0';
         else
            blk_lnk_up_d       <= blk_lnk_up; -- create delay of blk_lnk_up for edge detect
            if rdata_str_done_int = '1' then
               arid_rresp(cpl_index_int)      <= (others => '0');
            end if;
            if illegal_burst_int = '1' or bar_error_int = '1' then
               arid_rresp(rd_req_ptr)         <= "10"; -- SLVERR
            end if;
            if unsupported_req = '1' or completer_abort = '1' then
               arid_rresp(rd_req_index_err)   <= "10"; -- SLVERR
            end if;
            for i in 0 to C_AXIREAD_NUM-1 loop
               if cpl_timer_timeout_strb_int(i) = '1' or poisoned_req(i) = '1' or
                  (blk_lnk_up = '0' and blk_lnk_up_d = '1' and
                  not(i = cpl_index_int and en_rresp = '1' and read_dataSM_cs_d = STR_DATA)
                  and ((pending_rd_reqs(i) = '1' and not(i = cpl_index_int and (rdata_str_done_int = '1' or clr_pending_rd_reqs_entry = '1')))
                       or (i = rd_req_ptr and en_barhit = '1')))
                  then --falling edge of blk_lnk_up, set if not current rresp
                  arid_rresp(i)                  <= "10"; -- SLVERR
               end if;
               if pending_rd_reqs(i) = '1' and pending_rd_reqs_d(i) = '0' and blk_lnk_up = '0' then --pending read req set during link down
                  arid_rresp(i)                  <= "10"; -- SLVERR
               end if;
            end loop;
         end if;
      end if;
   end process;

   -- This process maintains completion permission status for each 'slot' read request
   -- As completion staus is cleared of any pending completions, the state of the master bridge write is checked and
   -- permission is granted if it is IDLE. If not, a request is made to the ordering logic. When a go comes back
   -- permission is then granted.
   completion_permission_proc :process(s_axi_aclk)
   variable index_save : integer range 0 to 8;
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            slave_cmpl_rdy_p            <= '0';
            cpl_req_index               <= 0;
            cpl_permit                  <= (others => '0');
            cmpl_rdy_pend               <= (others => '0');
            slave_cmpl_go_pend          <= '0';
         else
            slave_cmpl_rdy_p      <= '0';
            index_save := HISTORY_SIZE;
            for i in 0 to C_AXIREAD_NUM-1 loop
               if pending_rd_reqs_d(i) = '1' and ((tag_cpl_status_clr(i)(0 to DATA_SIZE*8-1) = ONES and tag_cpl_status_clr_d(i)(0 to DATA_SIZE*8-1) /= ONES)
               or blk_lnk_up = '0') and cpl_permit(i) = '0' then
                  index_save            := i;
               end if;
            end loop;
            if index_save /= HISTORY_SIZE then
               if master_wr_idle = '0' then
                  if slave_cmpl_go_pend = '0' and cmpl_rdy_pend = 0 then
                     slave_cmpl_rdy_p            <= '1';
                     slave_cmpl_go_pend          <= '1';
                     cpl_req_index               <= index_save;
                  else
                     cmpl_rdy_pend(index_save)   <= '1';
                  end if;
               else
                  cpl_permit(index_save)   <= '1';
               end if;
            end if; 
            index_save := HISTORY_SIZE;
            for i in 0 to C_AXIREAD_NUM-1 loop
               if cmpl_rdy_pend(i) = '1' then
                  index_save            := i;
               end if;
            end loop;
            if index_save /= HISTORY_SIZE then
               if master_wr_idle = '0' then
                  if slave_cmpl_go_pend = '0' then
                     slave_cmpl_rdy_p            <= '1';
                     slave_cmpl_go_pend          <= '1';
                     cpl_req_index               <= index_save;
                  end if;
               else
                  cpl_permit(index_save)      <= '1';
                  cmpl_rdy_pend(index_save)   <= '0';
               end if;
            end if;
            if slave_cmpl_go = '1' and slave_cmpl_go_pend = '1' then
               cpl_permit(cpl_req_index)   <= '1';
               cmpl_rdy_pend(cpl_req_index) <= '0';
               slave_cmpl_go_pend          <= '0';
            end if;
            if clr_pending_rd_reqs_entry = '1' then
               cpl_permit(cpl_index_int)   <= '0';
            end if;
            if illegal_burst_int = '1' or bar_error_int = '1' then
               cpl_permit(rd_req_ptr)      <= '1';--set so read return happens
            end if;
         end if;
      end if;
   end process;

   -- This process returns the read data requested to the AXI read data channel
   -- Works with both the 'sync' and 'rd_counter' processes below 
   read_dataSM_comb :process(read_dataSM_cs, rdata, s_axi_rready, rd_counter, arlen_reg, cpl_index_int, slot_cleared,
                             pending_rd_reqs_d, tag_cpl_status_clr, arid_dependency, rdata_mask, poisoned_req,
                             clr_dependency_entry, new_dependency_entry, cpl_permit, master_wr_idle)
   variable first_zero : boolean;
   variable index_save : integer range 0 to HISTORY_SIZE;
   begin
      read_dataSM_ns        <= read_dataSM_cs;
      s_axi_rdata_int       <= (others => '0');
      s_axi_rlast_int       <= '0';
      en_rresp              <= '0';
      rvalid_int            <= '0';
      rdata_bram_rd_en_int  <= '0';
      rdata_str_done_int    <= '0';
      cpl_index_nxt         <= cpl_index_int;
      header_ep             <= '0';
      rdata_str_start       <= '0';
      ld_rd_counter         <= '0';
      case read_dataSM_cs is
         when IDLE =>
            if HISTORY_SIZE = 8 then
               if pending_rd_reqs_d /= x"00" then
                  read_dataSM_ns        <= WAIT_FOR_CPL;
               end if;
            else
               if pending_rd_reqs_d /= x"0" then
                  read_dataSM_ns        <= WAIT_FOR_CPL;
               end if;
            end if;

         when WAIT_FOR_CPL =>
            if clr_dependency_entry ='0' and new_dependency_entry = '0' then
               index_save := HISTORY_SIZE;
               first_zero := FALSE;
               for i in 0 to C_AXIREAD_NUM-1 loop
                  if pending_rd_reqs_d(i) = '1' and cpl_permit(i) = '1' and first_zero = FALSE and
                  arid_dependency(i) = HISTORY_SIZE then
                     index_save            := i;
                     first_zero            := TRUE;
                  end if;
               end loop;
               if index_save /= HISTORY_SIZE and master_wr_idle = '1' then
                  cpl_index_nxt         <= index_save;
                  read_dataSM_ns        <= LOAD_READ_COUNTER;
               end if;
            end if;
         when LOAD_READ_COUNTER =>
            ld_rd_counter         <= '1';
            read_dataSM_ns        <= FIRST_BRAM_READ;

         when FIRST_BRAM_READ =>
            rdata_str_start       <= '1';
            rdata_bram_rd_en_int  <= '1';
            read_dataSM_ns        <= STR_DATA;

         when STR_DATA =>
            rvalid_int            <= '1';
            en_rresp              <= '1';
            s_axi_rdata_int       <= rdata and rdata_mask;
            if rd_counter = 0 then
               s_axi_rlast_int       <= '1';
               if s_axi_rready = '1' then
                  read_dataSM_ns        <= STR_DONE;
                  if poisoned_req(cpl_index_int) = '1' then
                     header_ep             <= '1';
                  end if;
               end if;
            elsif s_axi_rready = '1' then
               rdata_bram_rd_en_int  <= '1';
            end if;

         when STR_DONE =>
            rdata_str_done_int    <= '1';
            read_dataSM_ns        <= WAIT_SLOT_CLR;

         when WAIT_SLOT_CLR =>
            if slot_cleared = '1' then
               read_dataSM_ns        <= IDLE;
            end if;

      end case;
   end process;

   -- This process returns the read data requested to the AXI read data channel
   -- Works with the 'comb' process above 
   read_dataSM_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            read_dataSM_cs        <= IDLE;
            read_dataSM_cs_d      <= IDLE;
            cpl_index_int         <= 0;
         else
            read_dataSM_cs        <= read_dataSM_ns;
            read_dataSM_cs_d      <= read_dataSM_cs;
            cpl_index_int         <= cpl_index_nxt;
         end if;
      end if;
   end process;

   rd_counter_proc : process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            rd_counter       <= 0;
         else
            if ld_rd_counter = '1' then
               rd_counter       <= conv_integer(arlen_reg(cpl_index_int)) + 1;
            elsif rdata_bram_rd_en_int = '1' then
               rd_counter       <= rd_counter - 1;
            end if;
         end if;
      end if;
   end process;

-- completion timer logic

-- change from v1_00_a, removes C_FAMILY test after spartan6 test
-- AXI ACLK @62.5Mhz case
cpl_timer_start_count <= 3125 when C_COMP_TIMEOUT = 0 and ((C_USER_CLK_FREQ = 1 and C_USER_CLK2_DIV2 = "FALSE") or (C_USER_CLK_FREQ = 2 and C_USER_CLK2_DIV2 = "TRUE")) else
                         3125000 when C_COMP_TIMEOUT = 1 and ((C_USER_CLK_FREQ = 1 and C_USER_CLK2_DIV2 = "FALSE") or (C_USER_CLK_FREQ = 2 and C_USER_CLK2_DIV2 = "TRUE")) else
-- AXI ACLK @125MHz case
--                         6250 when C_COMP_TIMEOUT = 0 else
-- Add in 2 us buffer (total of 250 clock cycles) 
-- (to account for GT latency on outgoing and incoming PCIe TLPs)
                         6500 when C_COMP_TIMEOUT = 0 else
                         6250000 when C_COMP_TIMEOUT = 1 else
                         0;

-- completion timers -- one for each AXI read request
   cpl_timers_rd_req : for j in 0 to C_AXIREAD_NUM-1 generate
      cpl_timers_str_size : for k in 0 to DATA_SIZE*8-1 generate


      cpl_timers_comb : process(cpl_timer_count(j,k), tag_cpl_status_clr(j)(k), tag_cpl_status_clr_d(j)(k), cpl_timer_start_count)
      begin
         cpl_timer_count_nxt(j,k)    <= cpl_timer_count(j,k);
         cpl_timer_timeout_int(j)(k)      <= '0';
         if tag_cpl_status_clr(j)(k) = '0' and tag_cpl_status_clr_d(j)(k) = '1' then
            cpl_timer_count_nxt(j,k)    <= cpl_timer_start_count;
         elsif cpl_timer_count(j,k) /= 0 and tag_cpl_status_clr(j)(k) = '0' then
            cpl_timer_count_nxt(j,k)    <= cpl_timer_count(j,k) - 1;
         elsif cpl_timer_count(j,k) = 0 and tag_cpl_status_clr(j)(k) = '0' then
            cpl_timer_timeout_int(j)(k)  <= '1';
         end if;
      end process;

      cpl_timers_sync : process(s_axi_aclk)
      begin
         if(rising_edge(s_axi_aclk)) then
            if(reset = '0') then
               cpl_timer_count(j,k)        <= 0;
               tag_cpl_status_clr_d(j)(k)   <= '0';
            else
               cpl_timer_count(j,k)        <= cpl_timer_count_nxt(j,k);
               tag_cpl_status_clr_d(j)(k)   <= tag_cpl_status_clr(j)(k);
            end if;
         end if;
      end process;

   end generate cpl_timers_str_size;
   end generate cpl_timers_rd_req;

   cpl_timer_timeout_delay : process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            cpl_timer_timeout_d       <= (others => '0');
         else
            cpl_timer_timeout_d       <= cpl_timer_timeout;
         end if;
      end if;
   end process;

   cpl_timer_timeout_strb_process : process(cpl_timer_timeout, cpl_timer_timeout_d)
   begin
      cpl_timer_timeout_strb_int    <= (others => '0');
      for j in 0 to C_AXIREAD_NUM-1 loop
         if cpl_timer_timeout(j) = '1' and cpl_timer_timeout_d(j) = '0' then
            cpl_timer_timeout_strb_int(j) <= '1';
         end if;
      end loop;
   end process;



end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_slave_write.vhd
--
-- Description:     
--                  
-- This VHDL file is the HDL design file for the AXI slave write bridge. 
--                   
--                  
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_slave_write.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.conv_std_logic_vector;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;


--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------



entity axi_slave_write is
   generic(
      --Family Generics
      C_FAMILY                : string  :="virtex7";
      C_S_AXI_ID_WIDTH        : integer := 4;
      C_S_AXI_ADDR_WIDTH      : integer := 32;
      C_S_AXI_DATA_WIDTH      : integer := 32;
      C_AXIBAR_NUM            : integer := 6;
      C_AXIBAR_0              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0     : std_logic_vector := x"0000_0000";
      C_AXIBAR_1              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1     : std_logic_vector := x"0000_0000";
      C_AXIBAR_2              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2     : std_logic_vector := x"0000_0000";
      C_AXIBAR_3              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3     : std_logic_vector := x"0000_0000";
      C_AXIBAR_4              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4     : std_logic_vector := x"0000_0000";
      C_AXIBAR_5              : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5     : std_logic_vector := x"0000_0000";
      C_AXIBAR_CHK_SLV_ERR    : string  := "FALSE"
   );
   port(

      -- AXI Global
      s_axi_aclk              : in  std_logic;
      reset                   : in  std_logic;

      -- AXI Slave Write Address Channel
      s_axi_awid              : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_awaddr            : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_awregion          : in  std_logic_vector(3 downto 0);
      s_axi_awlen             : in  std_logic_vector(7 downto 0);
      s_axi_awsize            : in  std_logic_vector(2 downto 0);
      s_axi_awburst           : in  std_logic_vector(1 downto 0);
      s_axi_awvalid           : in  std_logic;
      s_axi_awready           : out std_logic;

      -- AXI Slave Write Data Channel
      s_axi_wdata             : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_wstrb             : in  std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
      s_axi_wlast             : in  std_logic;
      s_axi_wvalid            : in  std_logic;
      s_axi_wready            : out std_logic;

      -- AXI Slave Write Response Channel
      s_axi_bid               : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_bresp             : out std_logic_vector(1 downto 0);
      s_axi_bvalid            : out std_logic;
      s_axi_bready            : in  std_logic;

      -- Ordering signals
      pend_slv_wr_cnt         : out std_logic_vector(1 downto 0);
      cmpl_slv_wr_cnt         : out std_logic_vector(1 downto 0);
      slv_write_idle          : out std_logic;
      -- internal interface
      wdata                   : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      wdata_valid             : out std_logic;
      first_word_offset       : out integer;
      wdata_fifo_full         : in  std_logic;
      wdata_fifo_allmost_full : in  std_logic;
      waddr                   : out std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      length_bytes            : out std_logic_vector(12 downto 0);
      wbarhit                 : out std_logic_vector(C_AXIBAR_NUM-1 downto 0);
      first_BE                : out std_logic_vector(3 downto 0);
      first_BE_valid          : out std_logic;
      last_BE                 : out std_logic_vector(3 downto 0);
      last_BE_valid           : out std_logic;
      wdata_str_done          : in  std_logic;
      wdata_str_start         : in  std_logic;
      illegal_burst           : out std_logic;
      illegal_burst_trns      : out std_logic;
      bar_error_trns          : out std_logic;
      block_trns_lnkdwn       : out std_logic;
      blk_lnk_up              : in  std_logic;
      m_axis_rw_tvalid        : in  std_logic;
      pcie_bme                : in  std_logic;
      tlp_str_start           : in  std_logic;  -- Indicates if Write Req TLP started to Enhanced bridge
      wr_ptr                  : out std_logic;
      rd_ptr                  : out std_logic
   );
end axi_slave_write;

architecture structure of axi_slave_write is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

   type addr_array_type is array (natural range <>) of std_logic_vector(31 downto 0);

   constant C_BAR_ADDR_MASK_ARRAY : addr_array_type := (
                             x"0000_0000" + C_AXIBAR_0 xnor C_AXIBAR_HIGHADDR_0, 
                             x"0000_0000" + C_AXIBAR_1 xnor C_AXIBAR_HIGHADDR_1, 
                             x"0000_0000" + C_AXIBAR_2 xnor C_AXIBAR_HIGHADDR_2, 
                             x"0000_0000" + C_AXIBAR_3 xnor C_AXIBAR_HIGHADDR_3, 
                             x"0000_0000" + C_AXIBAR_4 xnor C_AXIBAR_HIGHADDR_4, 
                             x"0000_0000" + C_AXIBAR_5 xnor C_AXIBAR_HIGHADDR_5);

   constant C_BAR_HIGHADDR_ARRAY : addr_array_type := (C_AXIBAR_HIGHADDR_0, 
                                                       C_AXIBAR_HIGHADDR_1, 
                                                       C_AXIBAR_HIGHADDR_2, 
                                                       C_AXIBAR_HIGHADDR_3, 
                                                       C_AXIBAR_HIGHADDR_4, 
                                                       C_AXIBAR_HIGHADDR_5);

   constant C_BAR_ARRAY : addr_array_type := (C_AXIBAR_0, 
                                              C_AXIBAR_1, 
                                              C_AXIBAR_2, 
                                              C_AXIBAR_3, 
                                              C_AXIBAR_4, 
                                              C_AXIBAR_5);

   type wid_array is array (0 to 1) of std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
   type waddr_array is array (0 to 1) of std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   type wregion_array is array (0 to 1) of std_logic_vector(3 downto 0);
   type wlength_array is array (0 to 1) of std_logic_vector(7 downto 0);
   type wsize_array is array (0 to 1) of std_logic_vector(2 downto 0);
   type wburst_array is array (0 to 1) of std_logic_vector(1 downto 0);
   type barhit_array is array (0 to 1) of std_logic_vector(C_AXIBAR_NUM-1 downto 0);

   signal wid_reg             : wid_array := ((others => '0'),(others => '0'));
   signal waddr_reg           : waddr_array;
   signal wregion_reg         : wregion_array;
   signal wlength_reg         : wlength_array;
   signal wsize_reg           : wsize_array;
   signal wburst_reg          : wburst_array;
   signal barhit_reg          : barhit_array;

   constant ZEROS             : std_logic_vector(5 downto 0) := "000000";
   signal barhit              : std_logic_vector(C_AXIBAR_NUM-1 downto 0);
   signal awready_int         : std_logic := '0';
   signal bvalid_ack          : std_logic := '0';
   signal en_bvalid           : std_logic;
   signal bvalid_int          : std_logic := '0';
   signal illegal_burst_int   : std_logic;
   signal illegal_burst_log   : std_logic_vector(1 downto 0);
   signal bar_error_int       : std_logic;
   signal bar_error_log       : std_logic_vector(1 downto 0);
   signal bresp_int           : wburst_array := ((others => '0'),(others => '0'));
   signal req_active          : std_logic;
   signal en_barhit           : std_logic;
   signal wr_req_ptr_in       : integer range 0 to 1 := 0;
   signal wr_req_ptr_out      : integer range 0 to 1 := 0;
   signal size                : integer range 1 to 16;
   signal num_beats           : integer range 1 to 16;
   signal beat_count          : integer range 0 to 16;
   signal en_first_wdata      : std_logic;
   signal en_wdata            : std_logic;
   signal write_done          : std_logic;

   constant NUM_STROBES       :integer := C_S_AXI_DATA_WIDTH/8;
   type strobe_array is array (0 to 3) of std_logic_vector(NUM_STROBES-1 downto 0);
   signal strobe_pipe         : strobe_array;
   --signal en_strobes0         : std_logic;
   --signal en_strobes1         : std_logic;
   signal en_strobes2         : std_logic;
   signal en_first_BE_valid   : std_logic;
   signal last_BE_valid_int   : std_logic;
   signal length_bytes_int        : std_logic_vector(12 downto 0);
   signal first_word_offset_int   : integer range 0 to (C_S_AXI_DATA_WIDTH/32-1) := 0; -- CR # 633509
   signal last_word_offset    : integer := 0; -- CR # 633509
   signal wdata_valid_int     : std_logic;
   signal en_wdata_d          : std_logic;
   signal s_axi_wready_int    : std_logic := '0';
   signal wr_req_ptr_in_inv   : integer range 0 to 1 := 0;
   signal wr_req_ptr_out_int  : integer range 0 to 1 := 0;
   signal blk_lnk_up_d        : std_logic;
   signal blk_lnk_down_reqs   : integer range 0 to 2;
   signal pend_slv_wr_cnt_int : std_logic_vector(1 downto 0);
   signal cmpl_slv_wr_cnt_int : std_logic_vector(1 downto 0);
   signal slv_write_idle_int  : std_logic;
   signal two_req_indicator   : std_logic;
   signal null_beat_count     : integer;
   signal address_offset      : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal find_first_word_offset : std_logic;

   signal wr_ptr_incr         : std_logic;
   signal rd_ptr_incr         : std_logic;
   signal normalize_rd_ptr    : std_logic;
   signal wr_ptr_int          : std_logic;
   signal rd_ptr_int          : std_logic;
   signal wdata_str_done_sticky : std_logic;
   signal wdata_str_start_sticky: std_logic;
   signal wdata_str_start_d   : std_logic;
   signal last_bresp_ok       : std_logic;
   signal wdata_str_done_and_bresp_ok : std_logic;

   -----------------------------------------------------------------------------
   -- State Machines
   -----------------------------------------------------------------------------

   type write_reqSM_STATES is (IDLE,
                               CHECK,
                               CHECK2,
                               ONE_REQ_ACTIVE,
                               TWO_REQ_ACTIVE);
   signal write_reqSM_cs : write_reqSM_STATES;
   signal write_reqSM_ns : write_reqSM_STATES;

   type first_BE_SM_STATES is (IDLE,
                               FIRST_BEAT);
   signal first_BE_SM_cs : first_BE_SM_STATES;
   signal first_BE_SM_ns : first_BE_SM_STATES;

   type write_dataSM_STATES is (IDLE,
                                FIRST_DATA_WORD,
                                DATA_STREAM,
                                DONE,
                                WAIT_TLP_START,
                                WAIT_STR_DONE,
                                FIRST_DATA_WORD_2,
                                DATA_STREAM_2,
                                DONE_2);
                                
   signal write_dataSM_cs : write_dataSM_STATES;
   signal write_dataSM_ns : write_dataSM_STATES;

-- This function calculates the number of ls byte enable bits that are zero
   function num_lsb_zeros(strobes : std_logic_vector(NUM_STROBES-1 downto 0))
                          return integer is
      variable count     : integer;
      variable first_one : boolean;
      variable i         : integer;
   begin
      first_one  := FALSE;
      count      := 0;
      for i in 0 to C_S_AXI_DATA_WIDTH/8-1 loop
         if (strobes(i) = '1'and (first_one = FALSE)) then
            first_one  := TRUE;
            count := 0 + i;
         end if;
         -- Nam - never hit condition -  we don't allow non-first data beat with no strobe
         -- NAM / JRH fixed typo. Was b 2.
         -- coverage off -item c 1 -condrow 2
         --if (not(first_one) and strobes(i) = '0') then
         --   count := count + 1;
         --end if;
      end loop;
      return(count);
   end function;

-- This function calculates the number of ms byte enable bits that are zero
   function num_msb_zeros(strobes : std_logic_vector(NUM_STROBES-1 downto 0))
                          return integer is
      variable count     : integer;
      variable first_one : boolean;
      variable i         : integer;
      constant LIMIT : integer := C_S_AXI_DATA_WIDTH/8;
   begin
      first_one  := FALSE;
      count      := LIMIT;
      for i in LIMIT-1 downto 0 loop
         if (strobes(i) = '1' and (first_one = FALSE)) then
            first_one  := TRUE;
            count := LIMIT - 1 - i;
         end if;
         -- Nam - never hit condition -  we don't allow non-first data beat with no strobe
         -- NAM / JRH fixed typo. Was b 2.
         -- coverage off -item c 1 -condrow 2
         --if (not(first_one) and strobes(i) = '0') then
            --count := count + 1;
         --end if;
      end loop;
      return(count);
   end function;


begin


   s_axi_awready          <= awready_int;
   s_axi_bvalid           <= bvalid_int;
   first_word_offset      <= first_word_offset_int;
   s_axi_bid              <= wid_reg(wr_req_ptr_out_int);
   wr_req_ptr_in_inv      <= 1 when wr_req_ptr_in = 0 else 0;
   s_axi_bresp            <= bresp_int(wr_req_ptr_out_int) when bvalid_ack = '1' and blk_lnk_up = '1' else
                             "10" when bvalid_ack = '1' and blk_lnk_up = '0' else -- SLVERR always when link down
                             (others => '0');

   length_bytes_int       <= SHL(("00000" & wlength_reg(wr_req_ptr_out)) + 1 - null_beat_count, conv_std_logic_vector(log2(C_S_AXI_DATA_WIDTH/8), 4))
                             - (first_word_offset_int + last_word_offset)*4;
   length_bytes           <= length_bytes_int;

   waddr                  <= address_offset(C_S_AXI_ADDR_WIDTH-1 downto 2) + waddr_reg(wr_req_ptr_out)(C_S_AXI_ADDR_WIDTH-1 downto 2) & "00"
                                when first_word_offset_int = 0
                             else address_offset(C_S_AXI_ADDR_WIDTH-1 downto 3) + waddr_reg(wr_req_ptr_out)(C_S_AXI_ADDR_WIDTH-1 downto 3) & "100"
                                when first_word_offset_int = 1
                             else address_offset(C_S_AXI_ADDR_WIDTH-1 downto 4) + waddr_reg(wr_req_ptr_out)(C_S_AXI_ADDR_WIDTH-1 downto 4) & "1000"
                                when first_word_offset_int = 2
                             else address_offset(C_S_AXI_ADDR_WIDTH-1 downto 4) + waddr_reg(wr_req_ptr_out)(C_S_AXI_ADDR_WIDTH-1 downto 4) & "1100";

   size                   <= C_S_AXI_DATA_WIDTH/8;
   num_beats              <= 1;
   last_BE_valid          <= last_BE_valid_int;-- when blk_lnk_up = '1' else '0';
   wbarhit                <= barhit_reg(wr_req_ptr_out);
   wdata_valid            <= wdata_valid_int;
   s_axi_wready           <= s_axi_wready_int;
   illegal_burst          <= illegal_burst_int;
   pend_slv_wr_cnt        <= pend_slv_wr_cnt_int;
   cmpl_slv_wr_cnt        <= cmpl_slv_wr_cnt_int;
   slv_write_idle         <= slv_write_idle_int;

   wr_ptr                 <= wr_ptr_int;
   rd_ptr                 <= rd_ptr_int;
   wdata_str_done_and_bresp_ok <= '1' when (wdata_str_done = '1' or wdata_str_done_sticky = '1') and (last_bresp_ok = '1') else '0';

   -- Get write address phase info from AXI for up to 2 "slots" when available
   -- Works with the 'sync' process below 
   write_reqSM_comb :process(write_reqSM_cs, s_axi_awvalid, wr_req_ptr_in, wr_req_ptr_out, s_axi_bready, bvalid_ack,
                             barhit, wburst_reg, blk_lnk_up, pcie_bme)
   begin
      write_reqSM_ns         <= write_reqSM_cs;
      awready_int            <= '0';
      req_active             <= '0';
      illegal_burst_int      <= '0';
      bar_error_int          <= '0';
      en_barhit              <= '0';
      slv_write_idle_int     <= '0';
      case write_reqSM_cs is

         when IDLE =>
            slv_write_idle_int     <= '1';
            if blk_lnk_up = '1' and pcie_bme = '1' then -- only assert awready if link is up
               awready_int            <= '1';
            end if;
            if s_axi_awvalid = '1' and blk_lnk_up = '1' and pcie_bme = '1' then
               -- aquire write req qualifiers
               write_reqSM_ns         <= CHECK;
               slv_write_idle_int     <= '0';
            end if;

         when CHECK =>
            -- check qualifiers
            en_barhit              <= '1';
            -- coverage off
            -- never hit, remove in 13.3
            if barhit = ZEROS(C_AXIBAR_NUM - 1 downto 0) then
               if (C_AXIBAR_CHK_SLV_ERR = "TRUE") then
                  bar_error_int          <= '1';
                  write_reqSM_ns         <= ONE_REQ_ACTIVE;
               else
                  bar_error_int          <= '0';
                  write_reqSM_ns         <= IDLE;
               end if;
            else
            -- coverage on
               write_reqSM_ns         <= ONE_REQ_ACTIVE;
            end if;
            if (wburst_reg(wr_req_ptr_in) /= "01") then
               illegal_burst_int      <= '1';
            end if;

         when CHECK2 =>
            -- check qualifiers
            en_barhit              <= '1';
            -- coverage off
            -- never hit, remove in 13.3
            if barhit = ZEROS(C_AXIBAR_NUM - 1 downto 0) then
               if (C_AXIBAR_CHK_SLV_ERR = "TRUE") then
                  bar_error_int     <= '1';
                  if bvalid_ack = '1' then
                     write_reqSM_ns <= ONE_REQ_ACTIVE;
                  else
                     write_reqSM_ns <= TWO_REQ_ACTIVE;
                  end if;
               else
                  bar_error_int  <= '0';
                  write_reqSM_ns <= ONE_REQ_ACTIVE;
               end if;
            -- coverage on
            elsif bvalid_ack = '1' then
               write_reqSM_ns <= ONE_REQ_ACTIVE;
            else
               write_reqSM_ns <= TWO_REQ_ACTIVE;
            end if;
            
            if (wburst_reg(wr_req_ptr_in) /= "01") then
               illegal_burst_int      <= '1';
            end if;

         when ONE_REQ_ACTIVE =>
            req_active             <= '1';
            if blk_lnk_up = '1' and pcie_bme = '1' then -- only assert awready if link is up
               awready_int            <= '1';
            end if;
            if s_axi_awvalid = '1' and blk_lnk_up = '1' and pcie_bme = '1' then
               -- aquire write req qualifiers
               if bvalid_ack = '0' then
                  write_reqSM_ns <= CHECK2;
               else
                  write_reqSM_ns <= CHECK;
               end if;
            elsif bvalid_ack = '1' then
               write_reqSM_ns <= IDLE;
            end if;

         when TWO_REQ_ACTIVE =>
            req_active <= '1';
            if bvalid_ack = '1' then
               write_reqSM_ns <= ONE_REQ_ACTIVE;
            end if;

      end case;
   end process;

   -- Get write address phase info from AXI for up to 2 "slots" when available
   -- Works with the 'comb' process above 
   write_reqSM_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            write_reqSM_cs        <= IDLE;
            wr_req_ptr_in         <= 0;
            wr_req_ptr_out        <= 0;
            wr_req_ptr_out_int    <= 0;
            wid_reg               <= (others => (others => '0'));
            waddr_reg             <= (others => (others => '0'));
            wregion_reg           <= (others => (others => '0'));
            wlength_reg           <= (others => (others => '0'));
            wsize_reg             <= (others => (others => '0'));
            wburst_reg            <= (others => (others => '0'));
            barhit_reg            <= (others => (others => '0'));
         else
            write_reqSM_cs <= write_reqSM_ns;
            if s_axi_awvalid = '1' and awready_int = '1' then
               wid_reg(wr_req_ptr_in)      <= s_axi_awid;
               waddr_reg(wr_req_ptr_in)    <= s_axi_awaddr;
               wregion_reg(wr_req_ptr_in)  <= s_axi_awregion;
               wlength_reg(wr_req_ptr_in)  <= s_axi_awlen;
               wsize_reg(wr_req_ptr_in)    <= s_axi_awsize;
               wburst_reg(wr_req_ptr_in)   <= s_axi_awburst;
            end if;
            
            if tlp_str_start = '1' then
               if wr_req_ptr_out = 0 then
                  wr_req_ptr_out        <= 1;
               else
                  wr_req_ptr_out        <= 0;
               end if;
            end if;
            if bvalid_ack = '1' then
               if wr_req_ptr_out_int = 0 then
                  wr_req_ptr_out_int   <= 1;
               else
                  wr_req_ptr_out_int   <= 0;
               end if;
            end if;
            if en_barhit = '1' then
               barhit_reg(wr_req_ptr_in)   <= barhit;
               if wr_req_ptr_in = 0 then
                  wr_req_ptr_in         <= 1;
               else
                  wr_req_ptr_in         <= 0;
               end if;
            end if;
         end if;
      end if;
   end process;

   two_req_indicator_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if reset = '0' or ((write_reqSM_cs = CHECK2 or write_reqSM_cs = TWO_REQ_ACTIVE) and bvalid_ack = '1') then
            two_req_indicator      <= '0';
         elsif write_reqSM_cs = ONE_REQ_ACTIVE and s_axi_awvalid = '1' and blk_lnk_up = '1' and pcie_bme = '1' and bvalid_ack = '0' then
            two_req_indicator      <= '1';
         end if;
      end if;
   end process;


   BAR_decoder :process(waddr_reg, wr_req_ptr_in)
--   Remove the use of AwRegion
--   BAR_decoder :process(wregion_reg, wr_req_ptr_in)
--   variable region    : integer;
--   begin
--      region                 := conv_integer(wregion_reg(wr_req_ptr_in));
--      barhit                 <= (others => '0');
--      -- Nam - always true if statement below
--      -- NAM / JRH fixed typo. Was b 2.
--      -- coverage off -item b 1 -allfalse
--      if region < C_AXIBAR_NUM then
--         barhit(region)         <= '1';
--      end if;
   variable address : integer;
   begin
--     address := conv_integer(waddr_reg(wr_req_ptr_in));
     barhit <= (others => '0');

     -- Nam - always true if statement below
     -- NAM /JRH fixed typo. Was b 2.
     -- coverage off -item b 1 -allfalse
     for i in 0 to (C_AXIBAR_NUM-1) loop
       if((waddr_reg(wr_req_ptr_in) <= C_BAR_HIGHADDR_ARRAY(i)) and (waddr_reg(wr_req_ptr_in) >= C_BAR_ARRAY(i))) then
         barhit(i) <= '1';
       end if;
     end loop;       
      
   end process;

   -- Make sure that write with an illegal burst or misses BAR does not generate MemWr TLP(s)
   -- Also do not generate MemWr TLP(s)for writes in process when link goes down
   illegal_burst_proccess : process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            illegal_burst_log                    <= (others => '0');
            bar_error_log                        <= (others => '0');
            blk_lnk_up_d                         <= '0';
            blk_lnk_down_reqs                    <= 0;
         else
            blk_lnk_up_d                         <= blk_lnk_up;
            if (C_AXIBAR_CHK_SLV_ERR = "TRUE") then
               if(illegal_burst_int = '1') then
                  illegal_burst_log(wr_req_ptr_in)     <= '1';
               end if;
               if(bar_error_int = '1') then
                  bar_error_log(wr_req_ptr_in)         <= '1';
               end if;
               if bvalid_ack = '1' then
                  illegal_burst_log(wr_req_ptr_out_int)<= '0';
                  bar_error_log(wr_req_ptr_out_int)    <= '0';
               end if;
            else
               if(illegal_burst_int = '1') then
                  illegal_burst_log(wr_req_ptr_in)     <= '1';
               
               elsif bvalid_ack = '1' then
                  illegal_burst_log(wr_req_ptr_out_int)<= '0';
               end if;
            end if;
            if blk_lnk_up_d = '1' and blk_lnk_up = '0' then
               if slv_write_idle_int = '0' then
                  if two_req_indicator = '1' and bvalid_ack = '0' then
                     blk_lnk_down_reqs                    <= 2;
                  elsif two_req_indicator = '1' then
                     blk_lnk_down_reqs                    <= 1;
                  elsif bvalid_ack = '0' then
                     blk_lnk_down_reqs                    <= 1;
                  else
                     blk_lnk_down_reqs                    <= 0;
                  end if;
               else
                  blk_lnk_down_reqs                    <= 0;
               end if;
            end if;
            if bvalid_ack = '1' and blk_lnk_down_reqs /= 0 then
               blk_lnk_down_reqs                    <= blk_lnk_down_reqs-1;
            end if;
         end if;
      end if;
   end process;

   block_trns_lnkdwn <= '1' when blk_lnk_down_reqs /=0 else '0';

   illegal_burst_trns     <= illegal_burst_log(wr_req_ptr_out);
   bar_error_trns         <= bar_error_log(wr_req_ptr_out);

   bresp_gen :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            bresp_int          <= (others => (others => '0')); -- OKAY is default
         else
            if bvalid_ack = '1' then -- clear bresp after assertion
               bresp_int(wr_req_ptr_out_int)  <= "00"; -- OKAY
            end if;
            if illegal_burst_int = '1' or bar_error_int = '1' then
               bresp_int(wr_req_ptr_in)       <= "10"; -- SLVERR
            end if;
            if blk_lnk_up_d = '1' and blk_lnk_up = '0' and slv_write_idle_int = '0' then
               if two_req_indicator = '1' and bvalid_ack = '0' then
                  bresp_int                      <= (others => "10"); -- SLVERR on both
               elsif two_req_indicator = '1' then
                  if wr_req_ptr_out_int = 0 then
                     bresp_int(1)          <= "10"; -- SLVERR on one active
                  else
                     bresp_int(0)          <= "10"; -- SLVERR on one active
                  end if;
               elsif bvalid_ack = '0' then
                  bresp_int(wr_req_ptr_out_int) <= "10"; -- SLVERR on one active
               end if;
            end if;
         end if;
      end if;
   end process;

   -- This process gets the write data from the AXI write data channel and enables writing into the Write FIFO
   -- Works with the 'sync' process below 
   write_dataSM_comb :process(  write_dataSM_cs, req_active, s_axi_wvalid, 
                   s_axi_wlast, s_axi_bready,
                                wdata_fifo_full, wdata_str_start, 
                                tlp_str_start, two_req_indicator, 
                                bvalid_ack, en_bvalid, 
                                wdata_str_done_and_bresp_ok, wdata_str_start_sticky,
                                last_bresp_ok)
   begin
      write_dataSM_ns       <= write_dataSM_cs;
      s_axi_wready_int      <= '0';
      en_first_wdata        <= '0';
      en_wdata              <= '0';
      write_done            <= '0';
      en_bvalid             <= '0';
      rd_ptr_incr           <= '0';
      wr_ptr_incr           <= '0';
      normalize_rd_ptr      <= '0';

      -- Assert BVALID once 1st Beat of Last splitted write TLP or 
      -- write TLP( in case of no split) is presented on AXI-S RW interface
      if (wdata_str_start = '1' or wdata_str_start_sticky = '1') and 
         (bvalid_ack = '0' and last_bresp_ok = '0') then
        en_bvalid <= '1';
      end if;

      case write_dataSM_cs is

         when IDLE =>
         
            -- Only check req_active in IDLE state
            if req_active = '1' then
               write_dataSM_ns    <= FIRST_DATA_WORD;
            end if;

         when FIRST_DATA_WORD =>

            s_axi_wready_int          <= '1';
            if s_axi_wvalid = '1' then
               en_first_wdata         <= '1';
               if s_axi_wlast = '1' then
                  write_dataSM_ns     <= DONE;
               else
                  write_dataSM_ns     <= DATA_STREAM;
               end if;
            end if;

         when DATA_STREAM =>

               s_axi_wready_int       <= '1';
               if s_axi_wvalid = '1' then
                  en_wdata            <= '1';
                  
                  -- If last beat then go to DONE,
                  -- otherwise stay in this state to capture data.
                  if s_axi_wlast = '1' then
                     write_dataSM_ns  <= DONE;
                  end if;
               end if;

         -- Done capturing data from AXI
         when DONE =>

            write_done <= '1';
            write_dataSM_ns <= WAIT_TLP_START;

         -- Wait for Enhanced TLP logic to start processing data stream.
         when WAIT_TLP_START =>
         
            -- Wait for indicator that TLP SM has recognized the TLP
            -- packet to start sending it to the Enhanced Bridge.
            if tlp_str_start = '1' then

               -- If more than 1 write request,
               -- start the process of capturing write data of 2nd request
               -- in another buffer else go to WAIT_STR_DONE state
               if two_req_indicator = '1' then
                  write_dataSM_ns <= FIRST_DATA_WORD_2;
               else
                  write_dataSM_ns <= WAIT_STR_DONE;
               end if;
            end if;

         -- In this state waiting for Enhanced Bridge to complete stream.
         -- However, if we see a new request, buffer in the data.
         when WAIT_STR_DONE =>
            
            -- Change priority here.
            -- If TLP data phase completes, go back to IDLE/FIRST_DATA_WORD
            -- based on req_active
            if wdata_str_done_and_bresp_ok = '1' then

               normalize_rd_ptr <= '1';

               -- Either no pending transfers
               -- or req_active is HIGH which might go LOW or remain HIGH on next cycle
               -- Go to IDLE in any case
               write_dataSM_ns <= IDLE;
            
            -- if we see a new request, buffer in the data of new request in another buffer
            elsif two_req_indicator = '1' then
                write_dataSM_ns <= FIRST_DATA_WORD_2;
            end if;
            
         -- See next address write to send to Enhanced Bridge
         -- Only get to this state if subsequent write to process.
         when FIRST_DATA_WORD_2 =>
           
            -- See if prior write request completes then go back to FIRST_DATA_WORD
            if wdata_str_done_and_bresp_ok = '1' then
               
               write_dataSM_ns <= FIRST_DATA_WORD;
               normalize_rd_ptr <= '1';
               
            else
               s_axi_wready_int <= '1';
               if s_axi_wvalid = '1' then
                  en_first_wdata   <= '1';
                  wr_ptr_incr      <= '1';
                  if s_axi_wlast = '1' then
                     write_dataSM_ns  <= DONE_2;
                  else
                     write_dataSM_ns  <= DATA_STREAM_2;
                  end if;
               end if;
            end if;

         -- Capturing 2nd data stream from AXI
         when DATA_STREAM_2 =>

               s_axi_wready_int <= '1';
               if s_axi_wvalid = '1' then
                  en_wdata <= '1';
                  
                  -- If we see the WLAST on the 2nd AXI write stream.
                  if s_axi_wlast = '1' then
                     write_dataSM_ns  <= DONE_2;
                  end if;
               end if;

         -- Done accepting 2nd AXI write data stream.
         when DONE_2 =>

            -- write_done flag must be high when we are done with streaming out MWr TLP(s) in full
            -- along with the response back for the earlier TLP.
            if wdata_str_done_and_bresp_ok = '1' then
               write_done  <= '1';
               write_dataSM_ns <= WAIT_TLP_START;
               rd_ptr_incr <= '1';
            end if;

         -- Default state
         when others =>

            write_dataSM_ns <= IDLE;

      end case;
   end process;

   -- This process gets the write data from the AXI write data channel and enables writing into the Write FIFO
   -- Works with the 'comb' process above 
   write_dataSM_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            write_dataSM_cs          <= IDLE;
            wdata_str_start_sticky   <= '0';
            wdata_str_start_d        <= '0';
            wdata_str_done_sticky    <= '0';
            last_bresp_ok            <= '0';
            rd_ptr_int               <= '0';
            wr_ptr_int               <= '0';
            bvalid_ack               <= '0';
            bvalid_int               <= '0';
         else
            write_dataSM_cs          <= write_dataSM_ns;
            wdata_str_start_d        <= wdata_str_start;
            
            -- Detect the posedge of wdata_str_start and maintain wdata_str_start_sticky HIGH
            -- till we get bvalid_ack back.
            if bvalid_ack = '1' then
               wdata_str_start_sticky <= '0';
            elsif wdata_str_start = '1' and wdata_str_start_d = '0' then
               wdata_str_start_sticky <= '1';
            end if;

            -- wdata_str_done is a single cycle pulse,
            -- register this signal and make it sticky in the sense that it will
            -- de-assert only when response is given back to AXI side 
            if wdata_str_done = '1' then
               wdata_str_done_sticky <= '1';
            end if;
           
            -- Assert last_bresp_ok when response is given back for any write request
            if bvalid_int = '1' and s_axi_bready = '1' then
               last_bresp_ok         <= '1';
            end if;
            
            if write_dataSM_cs = WAIT_TLP_START or write_dataSM_cs = IDLE then
               wdata_str_done_sticky <= '0';
               last_bresp_ok         <= '0';
            end if;
            
            -- Toggle rd_ptr_int if rd_ptr_incr is HIGH
            if rd_ptr_incr = '1' then
               if rd_ptr_int = '1' then
                  rd_ptr_int         <= '0';
               else
                  rd_ptr_int         <= '1';
               end if;
            end if;

            -- Toggle wr_ptr_int if wr_ptr_incr is HIGH
            if wr_ptr_incr = '1' then
               if wr_ptr_int = '1' then
                  wr_ptr_int         <= '0';
               else
                  wr_ptr_int         <= '1';
               end if;
            end if;

            -- Normalize rd_ptr_int
            if normalize_rd_ptr = '1' then
               rd_ptr_int            <= wr_ptr_int;
            end if;
            
            -- BVALID signal is acknowledged
            if en_bvalid = '1' and s_axi_bready = '1' then
               bvalid_ack            <= '1';
            else
               bvalid_ack            <= '0';
            end if;
           
            -- bvalid_int is an internal signal which is connected to s_axi_bvalid output
            if s_axi_bready = '1' and en_bvalid = '1' and bvalid_int = '1' then
               bvalid_int            <= '0';
            else
               bvalid_int            <= en_bvalid;
            end if;

         end if;
      end if;
   end process;


   -- Determine the value of first BE to be used in MemWr TLP generation
   -- Works with 'sync' process below
   first_BE_SM_comb :process(first_BE_SM_cs, en_first_wdata, en_wdata, size, beat_count, write_done, strobe_pipe(0))
   begin
      first_BE_SM_ns   <= first_BE_SM_cs;
      en_strobes2           <= '0';
      en_first_BE_valid     <= '0';
      case first_BE_SM_cs is
            when IDLE =>
               if en_first_wdata = '1' then
                  first_BE_SM_ns        <= FIRST_BEAT;
               end if;

            when FIRST_BEAT =>
               -- Wait until there's at least one valid data or it has reached end of data stream / zero length write
               if ( ( num_msb_zeros(strobe_pipe(0)) /= NUM_STROBES ) or ( write_done = '1' ) ) then
                  en_strobes2           <= '1';
                  first_BE_SM_ns        <= IDLE;
                  en_first_BE_valid     <= '1';
               end if;

      end case;
   end process;

   -- Determine the value of first BE to be used in MemWr TLP generation
   -- Works with 'comb' process above
   first_BE_SM_sync :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            first_BE_SM_cs        <= IDLE;
            first_BE              <= (others => '0');
            first_BE_valid        <= '0';
         else
            first_BE_SM_cs        <= first_BE_SM_ns;
            if en_first_wdata = '1' then
               first_BE              <= (others => '0');
            elsif en_strobes2 = '1' then
               if size = 4 then -- dword 32
                  first_BE <= strobe_pipe(0)(beat_count*4-1 downto beat_count*4-4);
               else -- 64/128
                  if num_lsb_zeros(strobe_pipe(0)) < 4 then
                     first_BE <= strobe_pipe(0)(3 downto 0);
                  elsif num_lsb_zeros(strobe_pipe(0)) < 8 and C_S_AXI_DATA_WIDTH >= 64 then
                     first_BE <= strobe_pipe(0)(7 downto 4);
                  elsif num_lsb_zeros(strobe_pipe(0)) < 12 and C_S_AXI_DATA_WIDTH = 128 then
                     first_BE <= strobe_pipe(0)(11 downto 8);
                  elsif C_S_AXI_DATA_WIDTH = 128 then
                     first_BE <= strobe_pipe(0)(15 downto 12);
                  end if;
               end if;
            end if;
            if en_first_BE_valid = '1' then
               first_BE_valid        <= '1';
            else
               first_BE_valid        <= '0';
            end if;
         end if;
      end if;
   end process;


   strobe_pipe_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0' or last_BE_valid_int = '1') then
            for i in 0 to 3 loop
               strobe_pipe(i)        <= (others => '0');
            end loop;
         elsif (en_first_wdata = '1' or en_wdata = '1') and num_msb_zeros(s_axi_wstrb) /= NUM_STROBES then
            strobe_pipe(0)        <= s_axi_wstrb;
            for i in 1 to 3 loop
               strobe_pipe(i)        <= strobe_pipe(i-1);
            end loop;
         end if;
      end if;
   end process;


   first_word_offset_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0' or last_BE_valid_int = '1') then
            first_word_offset_int     <= 0;
            find_first_word_offset    <= '0';
         elsif en_first_wdata = '1' or find_first_word_offset = '1' then
            if num_msb_zeros(s_axi_wstrb) = NUM_STROBES then -- null data beat case
               find_first_word_offset <= '1';
            else
               first_word_offset_int <= num_lsb_zeros(s_axi_wstrb)/4;
               find_first_word_offset <= '0';
            end if;
         end if;
      end if;
   end process;


   last_word_offset_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0' or last_BE_valid_int = '1') then
            last_word_offset     <= 0;
         elsif num_msb_zeros(s_axi_wstrb) = NUM_STROBES then -- null data beat case
            if num_msb_zeros(strobe_pipe(0)) = NUM_STROBES then
               last_word_offset  <= 0;
            else
               last_word_offset  <= num_msb_zeros(strobe_pipe(0))/4;
            end if;
         elsif s_axi_wlast = '1' and s_axi_wready_int = '1' then
            last_word_offset <= num_msb_zeros(s_axi_wstrb)/4;
         end if;
      end if;
   end process;

   -- Determine the value of last BE to be used in MemWr TLP generation, needs to have strobes from last write data beat
   last_BE_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            last_BE               <= (others => '0');
            last_BE_valid_int     <= '0';
         elsif write_done = '1' then
            if (en_first_BE_valid = '0') or (size > 4) then
               if size = 4 then -- dword 32
                  if length_bytes_int < 5 then -- 1 DW payload
                     last_BE            <= (others => '0');
                  else
                     last_BE            <= strobe_pipe(0)(beat_count*4-1 downto beat_count*4-4);
                  end if;
               elsif C_S_AXI_DATA_WIDTH >= 64 then -- 64/128
                  if num_msb_zeros(strobe_pipe(0)) < 4 then -- data in DW3
                     if num_lsb_zeros(strobe_pipe(0)) > NUM_STROBES-5 and length_bytes_int < 5 then
                        last_BE         <= (others => '0');
                     else
                        last_BE         <= strobe_pipe(0)(NUM_STROBES-1 downto NUM_STROBES-4);
                     end if;
                  elsif num_msb_zeros(strobe_pipe(0)) < 8 then -- data in DW2
                     if num_lsb_zeros(strobe_pipe(0)) > NUM_STROBES-9 and length_bytes_int < 5 then
                        last_BE         <= (others => '0');
                     else
                        last_BE         <= strobe_pipe(0)(NUM_STROBES-5 downto NUM_STROBES-8);
                     end if;
                  elsif C_S_AXI_DATA_WIDTH = 128 and num_msb_zeros(strobe_pipe(0)) < 12 then -- data in DW1
                     if num_lsb_zeros(strobe_pipe(0)) > NUM_STROBES-13 and length_bytes_int < 5 then
                        last_BE         <= (others => '0');
                     else
                        last_BE         <= strobe_pipe(0)(NUM_STROBES-9 downto NUM_STROBES-12);
                     end if;
                  elsif C_S_AXI_DATA_WIDTH = 128 then -- data in DW0
                     if length_bytes_int < 5 then
                        last_BE         <= (others => '0');
                     else
                        last_BE         <= strobe_pipe(0)(NUM_STROBES-13 downto NUM_STROBES-16);
                     end if;
                  end if;
               end if;
            else
               last_BE               <= (others => '0');
            end if;
            last_BE_valid_int     <= '1';
         else
            last_BE_valid_int     <= '0';
            last_BE               <= (others => '0');
         end if;
      end if;
   end process;


   write_databeat_counter :process(s_axi_aclk)
      variable temp_zeros : integer;
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            beat_count         <= 0;
            null_beat_count    <= 0;
         else
            temp_zeros            := num_lsb_zeros(s_axi_wstrb);
            if en_first_wdata = '1' then
               beat_count         <= 1;
               if num_msb_zeros(s_axi_wstrb) = NUM_STROBES then -- null data beat case
                  null_beat_count    <= 1;
               else
                  null_beat_count    <= 0;
               end if;
            elsif en_wdata = '1' then
               beat_count         <= 1;
               if num_msb_zeros(s_axi_wstrb) = NUM_STROBES then -- null data beat case
                  null_beat_count    <= null_beat_count + 1;
               end if;
            end if;
            if write_done = '1' then
               beat_count         <= 0;
            end if;
         end if;
      end if;
   end process;

   write_address_offset :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            address_offset     <= (others => '0');
         else
            if en_first_wdata = '1' then
               if num_msb_zeros(s_axi_wstrb) = NUM_STROBES then -- null data beat case
                  address_offset     <= conv_std_logic_vector(NUM_STROBES,C_S_AXI_ADDR_WIDTH);
               else
                  address_offset     <= (others => '0');
               end if;
            elsif en_wdata = '1' then
               if find_first_word_offset = '1' and num_msb_zeros(s_axi_wstrb) = NUM_STROBES then -- null data beat case
                  address_offset     <= address_offset + conv_std_logic_vector(NUM_STROBES,C_S_AXI_ADDR_WIDTH);
               end if;
            end if;
         end if;
      end if;
   end process;

   write_data_pipe :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            wdata           <= (others => '0');
         else
            if wdata_valid_int = '1' then
               wdata           <= (others => '0');
            end if;
            if en_wdata = '1' or en_first_wdata = '1' then
               for i in 0 to NUM_STROBES-1 loop
                  if s_axi_wstrb(i) = '1' then
                     wdata(i*8+7 downto i*8) <= s_axi_wdata(i*8+7 downto i*8);
                  end if;
               end loop;
            end if;
         end if;
      end if;
   end process;

   en_wdata_d_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            en_wdata_d      <= '0';
         elsif num_msb_zeros(s_axi_wstrb) /= NUM_STROBES then
            en_wdata_d      <= (en_wdata or en_first_wdata);
         else
            en_wdata_d      <= '0';
         end if;
      end if;
   end process;

   wdata_valid_int     <= en_wdata_d;

   -- Two 2-bit counters are maintained to indicate slave writes in process for the ordering logic
   -- When counts match, there are no writes in process
   ordering_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            pend_slv_wr_cnt_int      <= (others => '0');
            cmpl_slv_wr_cnt_int      <= (others => '0');
         else
            if s_axi_awvalid = '1' and awready_int = '1' then
               if pend_slv_wr_cnt_int = "11" then
                  pend_slv_wr_cnt_int      <= (others => '0');
               else
                  pend_slv_wr_cnt_int      <= pend_slv_wr_cnt_int + 1;
               end if;
            end if;
            if bvalid_ack = '1' then
               if cmpl_slv_wr_cnt_int = "11" then
                  cmpl_slv_wr_cnt_int      <= (others => '0');
               else
                  cmpl_slv_wr_cnt_int      <= cmpl_slv_wr_cnt_int + 1;
               end if;
            end if;
         end if;
      end if;
   end process;
end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        slave_bridge.vhd
--
-- Description:     
--                  
-- This VHDL file is the HDL design file for the AXI slave write bridge. 
--                   
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              slave_bridge.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.conv_integer;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;
use axi_pcie_v2_9_14.axi_pcie_mm_s_pkg.all;

library xpm;
use xpm.vcomponents.all;

entity slave_bridge is
   generic(
      --Family Generics
      C_FAMILY                      : string  :="virtex7";
      C_S_AXI_ID_WIDTH              : integer := 4;
      C_S_AXI_ADDR_WIDTH            : integer := 32;
      C_S_AXI_DATA_WIDTH            : integer := 32;
      C_M_AXIS_DATA_WIDTH           : integer := 32;
      C_COMP_TIMEOUT                : integer := 0; -- 0=50us, 1=50ms
      C_USER_CLK_FREQ               : integer := 1;
      C_USER_CLK2_DIV2              : string  := "FALSE";
      C_INCLUDE_RC                  : integer; -- := 0;
      C_S_AXI_SUPPORTS_NARROW_BURST : integer := 1;
      C_EP_LINK_PARTNER_RCB         : integer := 0;
      C_AXIREAD_NUM                 : integer := 8;  -- CR # 646225
      C_AXIBAR_NUM                  : integer := 6;
      C_AXIBAR_AS_0                 : integer := 0;
      C_AXIBAR_AS_1                 : integer := 0;
      C_AXIBAR_AS_2                 : integer := 0;
      C_AXIBAR_AS_3                 : integer := 0;
      C_AXIBAR_AS_4                 : integer := 0;
      C_AXIBAR_AS_5                 : integer := 0;
      C_AXIBAR_0                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0           : std_logic_vector := x"0000_0000";
      C_AXIBAR_1                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1           : std_logic_vector := x"0000_0000";
      C_AXIBAR_2                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2           : std_logic_vector := x"0000_0000";
      C_AXIBAR_3                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3           : std_logic_vector := x"0000_0000";
      C_AXIBAR_4                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4           : std_logic_vector := x"0000_0000";
      C_AXIBAR_5                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5           : std_logic_vector := x"0000_0000";
      C_AXIBAR_CHK_SLV_ERR          : string  := "FALSE"
   );
   port(

      -- AXI Global
      s_axi_aclk           : in  std_logic;
      reset                : in  std_logic;

      -- AXI Slave Write Address Channel
      s_axi_awid           : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_awaddr         : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_awregion       : in  std_logic_vector(3 downto 0);
      s_axi_awlen          : in  std_logic_vector(7 downto 0);
      s_axi_awsize         : in  std_logic_vector(2 downto 0);
      s_axi_awburst        : in  std_logic_vector(1 downto 0);
      s_axi_awvalid        : in  std_logic;
      s_axi_awready        : out std_logic;

      -- AXI Slave Write Data Channel
      s_axi_wdata          : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_wstrb          : in  std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
      s_axi_wlast          : in  std_logic;
      s_axi_wvalid         : in  std_logic;
      s_axi_wready         : out std_logic;

      -- AXI Slave Write Response Channel
      s_axi_bid            : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_bresp          : out std_logic_vector(1 downto 0);
      s_axi_bvalid         : out std_logic;
      s_axi_bready         : in  std_logic;

      -- AXI Slave Read Address Channel
      s_axi_arid           : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_araddr         : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_arregion       : in  std_logic_vector(3 downto 0);
      s_axi_arlen          : in  std_logic_vector(7 downto 0);
      s_axi_arsize         : in  std_logic_vector(2 downto 0);
      s_axi_arburst        : in  std_logic_vector(1 downto 0);
      s_axi_arvalid        : in  std_logic;
      s_axi_arready        : out std_logic;

      -- AXI Slave Read Data Channel
      s_axi_rid            : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_rdata          : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_rresp          : out std_logic_vector(1 downto 0);
      s_axi_rlast          : out std_logic;
      s_axi_rvalid         : out std_logic;
      s_axi_rready         : in  std_logic;

      -- AXIS Write Requester Channel
      m_axis_rw_tdata      : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_rw_tstrb      : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_rw_tlast      : out std_logic;
      m_axis_rw_tvalid     : out std_logic;
      m_axis_rw_tready     : in  std_logic;

      -- AXIS Read Requester Channel
      m_axis_rr_tid        : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      m_axis_rr_tdata      : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_rr_tstrb      : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_rr_tlast      : out std_logic;
      m_axis_rr_tvalid     : out std_logic;
      m_axis_rr_tready     : in  std_logic;

      -- AXIS Completion Requester Channel
      s_axis_rc_tdata      : in  std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      s_axis_rc_tstrb      : in  std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      s_axis_rc_tlast      : in  std_logic;
      s_axis_rc_tvalid     : in  std_logic;
      s_axis_rc_tready     : out std_logic;

      -- AXI2PCIE translation vectors
      axibar2pciebar0      : in  std_logic_vector(63 downto 0);
      axibar2pciebar1      : in  std_logic_vector(63 downto 0);
      axibar2pciebar2      : in  std_logic_vector(63 downto 0);
      axibar2pciebar3      : in  std_logic_vector(63 downto 0);
      axibar2pciebar4      : in  std_logic_vector(63 downto 0);
      axibar2pciebar5      : in  std_logic_vector(63 downto 0);

      -- AXI-S Block Interface
      blk_lnk_up           : in  std_logic;
      blk_bus_number       : in  std_logic_vector(7 downto 0);
      blk_device_number    : in  std_logic_vector(4 downto 0);
      blk_function_number  : in  std_logic_vector(2 downto 0);
      blk_command          : in  std_logic_vector(15 downto 0);
      blk_dcontrol         : in  std_logic_vector(15 downto 0);
      blk_lstatus          : in  std_logic_vector(15 downto 0);
      np_cpl_pending       : out std_logic;
      RP_bridge_en         : in  std_logic;

      -- Ordering signals
      --slrdready     : out std_logic;
      --slcplready     : out std_logic;
      --slrdsend             : in  std_logic;
      --slcplsend            : in  std_logic;
      pend_slv_wr_cnt      : out std_logic_vector(1 downto 0);
      cmpl_slv_wr_cnt      : out std_logic_vector(1 downto 0);
      wrreqpend            : in  std_logic_vector(2 downto 0);
      wrreqcomp            : in  std_logic_vector(2 downto 0);
      slv_write_idle       : out std_logic;
      s_axi_awvalid_o      : out std_logic;
      master_wr_idle       : in  std_logic;
      
      -- Interrupts
      SUR                  : out std_logic;
      SUC                  : out std_logic;
      SCT                  : out std_logic;
      SEP                  : out std_logic;
      SCA                  : out std_logic;
      SIB                  : out std_logic;
      config_gen_req       : in  std_logic
   );

end slave_bridge;

architecture structure of slave_bridge is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";


  component axi_pcie_v2_9_14_axi_upsizer
      generic(
          C_FAMILY                    : string  := "none";
          C_AXI_ID_WIDTH              : integer := 4;
          C_AXI_ADDR_WIDTH            : integer := 32;
          C_S_AXI_DATA_WIDTH          : integer := 32;
          C_M_AXI_DATA_WIDTH          : integer := 32;
          C_AXI_SUPPORTS_USER_SIGNALS : integer := 0;
          C_AXI_AWUSER_WIDTH          : integer := 1;
          C_AXI_ARUSER_WIDTH          : integer := 1;
          C_AXI_WUSER_WIDTH           : integer := 1;
          C_AXI_RUSER_WIDTH           : integer := 1;
          C_AXI_BUSER_WIDTH           : integer := 1;
          C_AXI_SUPPORTS_WRITE        : integer := 1;
          C_AXI_SUPPORTS_READ         : integer := 1;
          C_S_AXI_R_REGISTER        : integer := 0;        -- CR # 649227
          C_M_AXI_R_REGISTER        : integer := 0;        -- CR # 649227
          C_PACKING_LEVEL             : integer := 1;
          C_SUPPORT_BURSTS            : integer := 1;
          C_SINGLE_THREAD             : integer := 1
      );
      port(
     -- Globals
          ARESETN                     :in  std_logic;
          ACLK                        :in  std_logic;
     -- Slave Interface Write Address Ports
          S_AXI_AWID                  :in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          S_AXI_AWADDR                :in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
          S_AXI_AWLEN                 :in  std_logic_vector(7 downto 0);
          S_AXI_AWSIZE                :in  std_logic_vector(2 downto 0);
          S_AXI_AWBURST               :in  std_logic_vector(1 downto 0);
          S_AXI_AWLOCK                :in  std_logic_vector(1 downto 0);
          S_AXI_AWCACHE               :in  std_logic_vector(3 downto 0);
          S_AXI_AWPROT                :in  std_logic_vector(2 downto 0);
          S_AXI_AWREGION              :in  std_logic_vector(3 downto 0);
          S_AXI_AWQOS                 :in  std_logic_vector(3 downto 0);
          S_AXI_AWUSER                :in  std_logic_vector(0 downto 0);
          S_AXI_AWVALID               :in  std_logic;
          S_AXI_AWREADY               :out std_logic;
     -- Slave Interface Write Data Ports
          S_AXI_WDATA                 :in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
          S_AXI_WSTRB                 :in  std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
          S_AXI_WLAST                 :in  std_logic;
          S_AXI_WUSER                 :in  std_logic_vector(0 downto 0);
          S_AXI_WVALID                :in  std_logic;
          S_AXI_WREADY                :out std_logic;
     -- Slave Interface Write Response Ports
          S_AXI_BID                   :out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          S_AXI_BRESP                 :out std_logic_vector(1 downto 0);
          S_AXI_BUSER                 :out std_logic_vector(0 downto 0);
          S_AXI_BVALID                :out std_logic;
          S_AXI_BREADY                :in  std_logic;
     -- Slave Interface Read Address Ports
          S_AXI_ARID                  :in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          S_AXI_ARADDR                :in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
          S_AXI_ARLEN                 :in  std_logic_vector(7 downto 0);
          S_AXI_ARSIZE                :in  std_logic_vector(2 downto 0);
          S_AXI_ARBURST               :in  std_logic_vector(1 downto 0);
          S_AXI_ARLOCK                :in  std_logic_vector(1 downto 0);
          S_AXI_ARCACHE               :in  std_logic_vector(3 downto 0);
          S_AXI_ARPROT                :in  std_logic_vector(2 downto 0);
          S_AXI_ARREGION              :in  std_logic_vector(3 downto 0);
          S_AXI_ARQOS                 :in  std_logic_vector(3 downto 0);
          S_AXI_ARUSER                :in  std_logic_vector(0 downto 0);
          S_AXI_ARVALID               :in  std_logic;
          S_AXI_ARREADY               :out std_logic;
     -- Slave Interface Read Data Ports
          S_AXI_RID                   :out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          S_AXI_RDATA                 :out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
          S_AXI_RRESP                 :out std_logic_vector(1 downto 0);
          S_AXI_RLAST                 :out std_logic;
          S_AXI_RUSER                 :out std_logic_vector(0 downto 0);
          S_AXI_RVALID                :out std_logic;
          S_AXI_RREADY                :in  std_logic;
     -- Master Interface Write Address Port
          M_AXI_AWID                  :out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          M_AXI_AWADDR                :out std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
          M_AXI_AWLEN                 :out std_logic_vector(7 downto 0);
          M_AXI_AWSIZE                :out std_logic_vector(2 downto 0);
          M_AXI_AWBURST               :out std_logic_vector(1 downto 0);
          M_AXI_AWREGION              :out std_logic_vector(3 downto 0);
          M_AXI_AWUSER                :out std_logic_vector(0 downto 0);
          M_AXI_AWVALID               :out std_logic;
          M_AXI_AWREADY               :in  std_logic;
	  M_AXI_AWLOCK                :out std_logic_vector(1 downto 0);
	  M_AXI_AWCACHE               :out std_logic_vector(3 downto 0);
	  M_AXI_AWPROT                :out std_logic_vector(2 downto 0);
	  M_AXI_AWQOS                 :out std_logic_vector(3 downto 0);
     -- Master Interface Write Data Ports
          M_AXI_WDATA                 :out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
          M_AXI_WSTRB                 :out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0);
          M_AXI_WLAST                 :out std_logic;
          M_AXI_WUSER                 :out std_logic_vector(0 downto 0);
          M_AXI_WVALID                :out std_logic;
          M_AXI_WREADY                :in  std_logic;
     -- Master Interface Write Response Ports
          M_AXI_BID                   :in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          M_AXI_BRESP                 :in  std_logic_vector(1 downto 0);
          M_AXI_BUSER                 :in  std_logic_vector(0 downto 0);
          M_AXI_BVALID                :in  std_logic;
          M_AXI_BREADY                :out std_logic;
     -- Master Interface Read Address Port
          M_AXI_ARID                  :out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          M_AXI_ARADDR                :out std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
          M_AXI_ARLEN                 :out std_logic_vector(7 downto 0);
          M_AXI_ARSIZE                :out std_logic_vector(2 downto 0);
          M_AXI_ARBURST               :out std_logic_vector(1 downto 0);
          M_AXI_ARREGION              :out std_logic_vector(3 downto 0);
          M_AXI_ARUSER                :out std_logic_vector(3 downto 0);
          M_AXI_ARVALID               :out std_logic;
          M_AXI_ARREADY               :in  std_logic;
	  M_AXI_ARLOCK                :out std_logic_vector(1 downto 0);
	  M_AXI_ARCACHE               :out std_logic_vector(3 downto 0);
	  M_AXI_ARPROT                :out std_logic_vector(2 downto 0);
	  M_AXI_ARQOS                 :out std_logic_vector(3 downto 0);
     -- Master Interface Read Data Ports
          M_AXI_RID                   :in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
          M_AXI_RDATA                 :in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
          M_AXI_RRESP                 :in  std_logic_vector(1 downto 0);
          M_AXI_RLAST                 :in  std_logic;
          M_AXI_RUSER                 :in  std_logic_vector(0 downto 0);
          M_AXI_RVALID                :in  std_logic;
          M_AXI_RREADY                :out std_logic
     );
  end component;


-- CONSTANTS --

   constant RD_BUFFER_DEPTH         : integer := 256*C_AXIREAD_NUM; -- 4, 8 or 16 bytes wide
   constant RD_BUFFER_ADDR_SIZE     : integer := log2(RD_BUFFER_DEPTH);
   constant ONES                    : std_logic_vector(0 to C_S_AXI_DATA_WIDTH/4-1):= (others => '1');
   constant ZEROS                   : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0) := (others => '0');
   signal wdata_fifo_dout           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata_fifo_dout1          : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata_fifo_dout2          : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata_fifo_rd_en          : std_logic := '0'; 
   signal wdata_fifo_rd_en1         : std_logic := '0'; 
   signal wdata_fifo_rd_en2         : std_logic := '0'; 
   signal wdata_fifo_empty          : std_logic;
   signal wdata_fifo_empty1         : std_logic;
   signal wdata_fifo_empty2         : std_logic;
   signal wdata_fifo_almost_empty   : std_logic;
   signal wdata_fifo_full           : std_logic;
   signal wdata_fifo_full1          : std_logic;
   signal wdata_fifo_full2          : std_logic;
   signal wdata_fifo_allmost_full   : std_logic;
   signal wdata_fifo_allmost_full1  : std_logic;
   signal wdata_fifo_allmost_full2  : std_logic;

   signal wdata                     : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata1                    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata2                    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal wdata_valid               : std_logic;
   signal wdata_valid1              : std_logic;
   signal wdata_valid2              : std_logic;
   signal waddr                     : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal wlength_bytes             : std_logic_vector(12 downto 0);
   signal rlength_bytes             : std_logic_vector(12 downto 0);
   signal wbarhit                   : std_logic_vector(C_AXIBAR_NUM-1 downto 0);
   signal wfirst_BE                 : std_logic_vector(3 downto 0);
   signal wfirst_BE_valid           : std_logic;
   signal wlast_BE                  : std_logic_vector(3 downto 0);
   signal wlast_BE_valid            : std_logic;
   signal raddr                     : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal rbarhit                   : std_logic_vector(C_AXIBAR_NUM-1 downto 0);
   signal araddr_2lsbs              : std_logic_vector(1 downto 0);
   signal rlast_BE                  : std_logic_vector(3 downto 0);
   signal read_req_sent             : std_logic;
   signal tag_sent                  : std_logic_vector(7 downto 0);
   signal length_sent               : std_logic_vector(9 downto 0);
   signal rreq_active               : std_logic;
   signal req_active_ptr            : integer range 0 to C_AXIREAD_NUM-1;
   signal req_active_ptr_d          : integer range 0 to C_AXIREAD_NUM-1;
   signal rdata_bram_rd_en          : std_logic;
   signal rdata_bram_addr           : std_logic_vector(RD_BUFFER_ADDR_SIZE-1 downto 0);
   signal rdata                     : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal data_stream_out           : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
   signal cpl_buffer_addr           : std_logic_vector(RD_BUFFER_ADDR_SIZE-1 downto 0);
   signal cpl_data_str_done         : std_logic;
   signal tag_in_cpl                : std_logic_vector(7 downto 0);
   signal tag_cpl_status_clr        : tag_cpl_status_clr_array;
   signal tag_cpl_status_clr_d      : tag_cpl_status_clr_array;
   signal cpl_index                 : integer range 0 to C_AXIREAD_NUM-1;
   signal rdata_str_done            : std_logic;
   signal rdata_str_start           : std_logic;
   signal wdata_str_done            : std_logic;
   signal wdata_str_start           : std_logic;
   signal wfirst_word_offset        : integer;
   signal first_word_offset         : first_word_offset_array;
   signal reqID                     : std_logic_vector(15 downto 0) := x"5A5A";
   signal maxpayloadsize            : std_logic_vector(2 downto 0) := "000";
   signal maxreadreqsize            : std_logic_vector(2 downto 0) := "000";
   signal sig_m_axis_rr_tlast       : std_logic;
   signal wea                       : std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
   signal illegal_burst_wr          : std_logic;
   signal illegal_burst_rd          : std_logic;
   signal illegal_burst_trns_wr     : std_logic;
   signal illegal_burst_trns_rd     : std_logic;
   signal bar_error_rd              : std_logic;
   signal bar_error_trns_wr         : std_logic;
   signal bar_error_trns_rd         : std_logic;
   signal unsupported_req           : std_logic;
   signal unexpected_cpl            : std_logic;
   signal header_ep                 : std_logic;
   signal completer_abort           : std_logic;
   signal cpl_timer_timeout_strb    : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal rd_req_index_err          : integer range 0 to C_AXIREAD_NUM-1;
   signal poisoned_req              : std_logic_vector(C_AXIREAD_NUM-1 downto 0);
   signal reset_inv_wr_fifo         : std_logic;
   signal illegal_burst_int_wr      : std_logic;
   signal illegal_burst_int_rd      : std_logic;
   signal illegal_burst_int         : std_logic;
   signal block_trns_lnkdwn         : std_logic;

   -- Master Interface Write Address Port
   signal sig_m_axi_awid            : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
   signal sig_m_axi_awaddr          : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal sig_m_axi_awlen           : std_logic_vector(7 downto 0);
   signal sig_m_axi_awsize          : std_logic_vector(2 downto 0);
   signal sig_m_axi_awburst         : std_logic_vector(1 downto 0);
   signal sig_m_axi_awregion        : std_logic_vector(3 downto 0);
   signal sig_m_axi_awvalid         : std_logic;
   signal sig_m_axi_awready         : std_logic;
   -- Master Interface Write Data Ports
   signal sig_m_axi_wdata           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal sig_m_axi_wstrb           : std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
   signal sig_m_axi_wlast           : std_logic;
   signal sig_m_axi_wvalid          : std_logic;
   signal sig_m_axi_wready          : std_logic;
   -- Master Interface Write Response Ports
   signal sig_m_axi_bid             : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
   signal sig_m_axi_bresp           : std_logic_vector(1 downto 0);
   signal sig_m_axi_bvalid          : std_logic;
   signal sig_m_axi_bready          : std_logic;
   -- Master Interface Read Address Port
   signal sig_m_axi_arid            : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
   signal sig_m_axi_araddr          : std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
   signal sig_m_axi_arlen           : std_logic_vector(7 downto 0);
   signal sig_m_axi_arsize          : std_logic_vector(2 downto 0);
   signal sig_m_axi_arburst         : std_logic_vector(1 downto 0);
   signal sig_m_axi_arregion        : std_logic_vector(3 downto 0);
   signal sig_m_axi_arvalid         : std_logic;
   signal sig_m_axi_arready         : std_logic;
   -- Master Interface Read Data Ports
   signal sig_m_axi_rid             : std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
   signal sig_m_axi_rdata           : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
   signal sig_m_axi_rresp           : std_logic_vector(1 downto 0);
   signal sig_m_axi_rlast           : std_logic;  
   signal sig_m_axi_rvalid          : std_logic;
   signal sig_m_axi_rready          : std_logic;
   signal pend_slv_wr_cnt_sig         : std_logic_vector(1 downto 0);
   signal cmpl_slv_wr_cnt_sig         : std_logic_vector(1 downto 0);
   signal slrdreadycnt, slcplreadycnt : std_logic_vector(3 downto 0);
   signal slrdorderpipeline           : std_logic_vector(3 downto 0);
   signal slcplorderpipeline          : std_logic_vector(3 downto 0);
   signal slrdready, slcplready       : std_logic := '0';
   signal slrdsend, slcplsend         : std_logic;
   type mswrreqpendrecord_array is array (0 to 7) of std_logic_vector(2 downto 0);
   signal mswrreqpendrecord           : mswrreqpendrecord_array;
   type slwrreqpendrecord_array is array (0 to 7) of std_logic_vector(1 downto 0);
   signal slwrreqpendrecord           : slwrreqpendrecord_array;
   signal sig_slv_write_idle          : std_logic;
   signal sig_m_axis_rw_tvalid        : std_logic;
   signal total_length_out            : integer;
   signal tag_pending_for_cpl         : std_logic;
   signal tag_len_active_valid        : std_logic;
   signal sig_pcie_bme                : std_logic;
   signal sig_tlp_str_start           : std_logic;
   signal sig_m_axis_rr_tvalid        : std_logic;
   signal sig_np_cpl_pending          : std_logic_vector(0 to C_AXIREAD_NUM-1);
   signal wr_ptr                      : std_logic;
   signal rd_ptr                      : std_logic;
   signal pu_axi_arsize_d             : std_logic_vector(2 downto 0);
   signal pu_axi_arlen_d              : std_logic_vector(7 downto 0);
   signal sig_s_axi_arready           : std_logic;
   signal read_req_sent_array         : std_logic_vector(0 to C_AXIREAD_NUM-1);
   signal sig_SCT                     : std_logic;

begin

   m_axis_rr_tlast     <= sig_m_axis_rr_tlast;
   m_axis_rw_tvalid    <= sig_m_axis_rw_tvalid;
   m_axis_rr_tvalid    <= sig_m_axis_rr_tvalid;
   s_axi_awvalid_o     <= sig_m_axi_awvalid;
   reqID               <= blk_bus_number & blk_device_number & blk_function_number;
   maxpayloadsize      <= blk_dcontrol(7 downto 5);
   maxreadreqsize      <= blk_dcontrol(14 downto 12);
   reset_inv_wr_fifo   <= not(reset);

   pend_slv_wr_cnt     <= pend_slv_wr_cnt_sig;
   cmpl_slv_wr_cnt     <= cmpl_slv_wr_cnt_sig;
   slv_write_idle      <= sig_slv_write_idle;
   -- Interrupts
   SUR                 <= unsupported_req;
   SUC                 <= unexpected_cpl and reset;--block with reset
   SCT                 <= sig_SCT;
   SEP                 <= header_ep;
   SCA                 <= completer_abort;
   SIB                 <= illegal_burst_int;
   sig_pcie_bme        <= blk_command(2) when C_INCLUDE_RC = 0 else RP_bridge_en; --BME only if EP, use RP_bridge_en to block if RC

   np_cpl_pending      <= '0' when sig_np_cpl_pending = 0 else '1';

   -- wdata FIFO routing glue logic
   wdata1              <= wdata when wr_ptr = '0' else ZEROS;
   wdata2              <= wdata when wr_ptr = '1' else ZEROS;
   wdata_valid1        <= wdata_valid when wr_ptr = '0' else '0';
   wdata_valid2        <= wdata_valid when wr_ptr = '1' else '0';
   wdata_fifo_rd_en1   <= wdata_fifo_rd_en when rd_ptr = '0' else '0';
   wdata_fifo_rd_en2   <= wdata_fifo_rd_en when rd_ptr = '1' else '0';
   wdata_fifo_dout     <= wdata_fifo_dout1 when rd_ptr = '0' else wdata_fifo_dout2;
   wdata_fifo_allmost_full <= wdata_fifo_allmost_full1 when wr_ptr = '0' else wdata_fifo_allmost_full2;
   wdata_fifo_full     <= wdata_fifo_full1 when wr_ptr = '0' else wdata_fifo_full2;
   wdata_fifo_empty    <= wdata_fifo_empty1 when rd_ptr = '0' else wdata_fifo_empty2;

   np_cpl_pending_proc: process (s_axi_aclk)
   begin
      if rising_edge(s_axi_aclk) then
         if reset = '0' then
            sig_np_cpl_pending       <= (others => '0');
            tag_cpl_status_clr_d     <= (others => (others => '1'));
         else
            tag_cpl_status_clr_d     <= tag_cpl_status_clr;
            -- Set the slot in which request is registered
            --if sig_m_axis_rr_tvalid = '1' and m_axis_rr_tready = '1' then
            --   sig_np_cpl_pending(req_active_ptr) <= '1';
            --end if;
            -- Clear the slot for which request is completed
            for j in 0 to C_AXIREAD_NUM-1 loop
               if tag_cpl_status_clr(j)(0 to C_S_AXI_DATA_WIDTH/4-1) = ONES and 
                  tag_cpl_status_clr_d(j)(0 to C_S_AXI_DATA_WIDTH/4-1) /= ONES then 
                  sig_np_cpl_pending(j)  <= '0';
               end if;
            end loop;
            -- Set the slot in which request is registered
            if sig_m_axis_rr_tvalid = '1' and m_axis_rr_tready = '1' then
               sig_np_cpl_pending(req_active_ptr) <= '1';
            end if;
         end if;
      end if;
   end process;

   sct_proc: process (s_axi_aclk)
   begin
      if rising_edge(s_axi_aclk) then
         if reset = '0' then
            req_active_ptr_d    <= 0;
            read_req_sent_array <= (others => '0');
            sig_SCT             <= '0';
         else
            req_active_ptr_d    <= req_active_ptr;
            sig_SCT             <= '0';
            if read_req_sent = '1' then
               read_req_sent_array(req_active_ptr_d) <= '1';
            end if;
            if cpl_timer_timeout_strb /= 0 then
               for i in 0 to C_AXIREAD_NUM-1 loop
                  if cpl_timer_timeout_strb(i) = '1' and read_req_sent_array(i) = '1' then
                     sig_SCT <= '1';
                     read_req_sent_array(i) <= '0';
                  end if;
               end loop;
            end if;
         end if;
      end if;
   end process;

   slave_rd_ordering: process (s_axi_aclk)
   begin
      if rising_edge(s_axi_aclk) then
         if reset = '0' then
            slrdorderpipeline <= (others => '0');
            slrdsend <= '0';
            slrdreadycnt <= "0000";
         else
            if slrdready = '1' then
               slrdreadycnt <= slrdreadycnt + 1;
               slwrreqpendrecord(conv_integer(slrdreadycnt(2 downto 0))) <= pend_slv_wr_cnt_sig;
            end if;
            slrdsend <= '0';
            if slrdreadycnt /= slrdorderpipeline then
               if slwrreqpendrecord(conv_integer(slrdorderpipeline(2 downto 0))) = cmpl_slv_wr_cnt_sig then
                  slrdsend <= '1';
                  slrdorderpipeline <= slrdorderpipeline + 1;
               end if;
            end if;
         end if;
      end if;
   end process;

   slave_cpl_ordering: process (s_axi_aclk)
   begin
      if rising_edge(s_axi_aclk) then
         if reset = '0' then
            slcplorderpipeline <= (others => '0');
            slcplsend <= '0';
            slcplreadycnt <= "0000";
         else
            if slcplready = '1' then
               slcplreadycnt <= slcplreadycnt + 1;
               mswrreqpendrecord(conv_integer(slcplreadycnt(2 downto 0))) <= wrreqpend;
            end if;
            slcplsend <= '0';
            if slcplreadycnt /= slcplorderpipeline then
               if mswrreqpendrecord(conv_integer(slcplorderpipeline(2 downto 0))) = wrreqcomp then
                  slcplsend <= '1';
                  slcplorderpipeline <= slcplorderpipeline + 1;
               end if;
            end if;
         end if;
      end if;
   end process;

   illegal_burst_int_proc :process(s_axi_aclk)
   begin
      if(rising_edge(s_axi_aclk)) then
         if(reset = '0') then
            illegal_burst_int_wr     <= '0';
            illegal_burst_int_rd     <= '0';
            illegal_burst_int        <= '0';
         else
            if(illegal_burst_wr = '1') then
               illegal_burst_int_wr     <= '1';
            end if;
            if(illegal_burst_rd = '1') then
               illegal_burst_int_rd     <= '1';
            end if;
            if(illegal_burst_int_wr = '1' and illegal_burst_int = '0') then
               illegal_burst_int        <= '1';
               illegal_burst_int_wr     <= '0';
            elsif(illegal_burst_int_rd = '1' and illegal_burst_int = '0') then
               illegal_burst_int        <= '1';
               illegal_burst_int_rd     <= '0';
            else
               illegal_burst_int        <= '0';
            end if;
         end if;
      end if;
   end process;


   comp_axi_slave_write : entity axi_pcie_v2_9_14.axi_slave_write
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_S_AXI_ID_WIDTH        => C_S_AXI_ID_WIDTH,
      C_S_AXI_ADDR_WIDTH      => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH      => C_S_AXI_DATA_WIDTH,
      C_AXIBAR_NUM            => C_AXIBAR_NUM,
      C_AXIBAR_0              => C_AXIBAR_0,
      C_AXIBAR_HIGHADDR_0     => C_AXIBAR_HIGHADDR_0,
      C_AXIBAR_1              => C_AXIBAR_1,
      C_AXIBAR_HIGHADDR_1     => C_AXIBAR_HIGHADDR_1,
      C_AXIBAR_2              => C_AXIBAR_2,
      C_AXIBAR_HIGHADDR_2     => C_AXIBAR_HIGHADDR_2,
      C_AXIBAR_3              => C_AXIBAR_3,
      C_AXIBAR_HIGHADDR_3     => C_AXIBAR_HIGHADDR_3,
      C_AXIBAR_4              => C_AXIBAR_4,
      C_AXIBAR_HIGHADDR_4     => C_AXIBAR_HIGHADDR_4,
      C_AXIBAR_5              => C_AXIBAR_5,
      C_AXIBAR_HIGHADDR_5     => C_AXIBAR_HIGHADDR_5,
      C_AXIBAR_CHK_SLV_ERR    => C_AXIBAR_CHK_SLV_ERR
   )
   port map(

      -- AXI Global
      s_axi_aclk              => s_axi_aclk,
      reset                   => reset,

      -- AXI Slave Write Address Channel
      s_axi_awid              => sig_m_axi_awid,
      s_axi_awaddr            => sig_m_axi_awaddr,
      s_axi_awregion          => sig_m_axi_awregion,
      s_axi_awlen             => sig_m_axi_awlen,
      s_axi_awsize            => sig_m_axi_awsize,
      s_axi_awburst           => sig_m_axi_awburst,
      s_axi_awvalid           => sig_m_axi_awvalid,
      s_axi_awready           => sig_m_axi_awready,

      -- AXI Slave Write Data Channel
      s_axi_wdata             => sig_m_axi_wdata,
      s_axi_wstrb             => sig_m_axi_wstrb,
      s_axi_wlast             => sig_m_axi_wlast,
      s_axi_wvalid            => sig_m_axi_wvalid,
      s_axi_wready            => sig_m_axi_wready,

      -- AXI Slave Write Response Channel
      s_axi_bid               => sig_m_axi_bid,
      s_axi_bresp             => sig_m_axi_bresp,
      s_axi_bvalid            => sig_m_axi_bvalid,
      s_axi_bready            => sig_m_axi_bready,

      -- Ordering signals
      pend_slv_wr_cnt         => pend_slv_wr_cnt_sig,
      cmpl_slv_wr_cnt         => cmpl_slv_wr_cnt_sig,
      slv_write_idle          => sig_slv_write_idle,
      -- internal interface
      wdata                   => wdata,
      wdata_valid             => wdata_valid,
      first_word_offset       => wfirst_word_offset,
      wdata_fifo_full         => wdata_fifo_full,
      wdata_fifo_allmost_full => wdata_fifo_allmost_full,
      waddr                   => waddr,
      length_bytes            => wlength_bytes,
      wbarhit                 => wbarhit,
      first_BE                => wfirst_BE,
      first_BE_valid          => wfirst_BE_valid,
      last_BE                 => wlast_BE,
      last_BE_valid           => wlast_BE_valid,
      wdata_str_done          => wdata_str_done,
      wdata_str_start         => wdata_str_start,
      illegal_burst           => illegal_burst_wr,
      illegal_burst_trns      => illegal_burst_trns_wr,
      bar_error_trns          => bar_error_trns_wr,
      block_trns_lnkdwn       => block_trns_lnkdwn,
      blk_lnk_up              => blk_lnk_up,
      m_axis_rw_tvalid        => sig_m_axis_rw_tvalid,
      pcie_bme                => sig_pcie_bme,
      tlp_str_start           => sig_tlp_str_start,
      wr_ptr                  => wr_ptr,
      rd_ptr                  => rd_ptr
   );

   comp_axi_slave_read : entity axi_pcie_v2_9_14.axi_slave_read
   generic map(
      --Family Generics
      C_FAMILY                      => C_FAMILY,
      C_S_AXI_ID_WIDTH              => C_S_AXI_ID_WIDTH,
      C_S_AXI_ADDR_WIDTH            => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH            => C_S_AXI_DATA_WIDTH,
      C_COMP_TIMEOUT                => C_COMP_TIMEOUT,
      C_USER_CLK_FREQ               => C_USER_CLK_FREQ,
      C_USER_CLK2_DIV2              => C_USER_CLK2_DIV2,
      C_S_AXI_SUPPORTS_NARROW_BURST => C_S_AXI_SUPPORTS_NARROW_BURST,
      C_AXIREAD_NUM                 => C_AXIREAD_NUM,
      C_RD_BUFFER_ADDR_SIZE         => RD_BUFFER_ADDR_SIZE,
      C_AXIBAR_NUM                  => C_AXIBAR_NUM,
      C_AXIBAR_0                    => C_AXIBAR_0,
      C_AXIBAR_HIGHADDR_0           => C_AXIBAR_HIGHADDR_0,
      C_AXIBAR_1                    => C_AXIBAR_1,
      C_AXIBAR_HIGHADDR_1           => C_AXIBAR_HIGHADDR_1,
      C_AXIBAR_2                    => C_AXIBAR_2,
      C_AXIBAR_HIGHADDR_2           => C_AXIBAR_HIGHADDR_2,
      C_AXIBAR_3                    => C_AXIBAR_3,
      C_AXIBAR_HIGHADDR_3           => C_AXIBAR_HIGHADDR_3,
      C_AXIBAR_4                    => C_AXIBAR_4,
      C_AXIBAR_HIGHADDR_4           => C_AXIBAR_HIGHADDR_4,
      C_AXIBAR_5                    => C_AXIBAR_5,
      C_AXIBAR_HIGHADDR_5           => C_AXIBAR_HIGHADDR_5,
      C_AXIBAR_CHK_SLV_ERR          => C_AXIBAR_CHK_SLV_ERR
   )
   port map(
      -- AXI Global
      s_axi_aclk              => s_axi_aclk,
      reset                   => reset,

      -- AXI Slave Read Address Channel
      s_axi_arid              => sig_m_axi_arid,
      s_axi_araddr            => sig_m_axi_araddr,
      s_axi_arregion          => sig_m_axi_arregion,
      s_axi_arlen             => sig_m_axi_arlen,
      s_axi_arsize            => sig_m_axi_arsize,
      s_axi_arburst           => sig_m_axi_arburst,
      s_axi_arvalid           => sig_m_axi_arvalid,
      s_axi_arready           => sig_m_axi_arready,
      pu_axi_arlen            => pu_axi_arlen_d,
      pu_axi_arsize           => pu_axi_arsize_d,

      -- AXI Slave Read Data Channel
      s_axi_rid               => sig_m_axi_rid,
      s_axi_rdata             => sig_m_axi_rdata,
      s_axi_rresp             => sig_m_axi_rresp,
      s_axi_rlast             => sig_m_axi_rlast,
      s_axi_rvalid            => sig_m_axi_rvalid,
      s_axi_rready            => sig_m_axi_rready,
      -- AXIS Read Requester Channel
      m_axis_rr_tid           => m_axis_rr_tid,
      -- Ordering signals
      slave_read_req_p        => slrdready,
      slave_rd_req_go         => slrdsend,
      slave_cmpl_rdy_p        => slcplready,
      slave_cmpl_go           => slcplsend,
      slv_write_idle          => sig_slv_write_idle,
      master_wr_idle          => master_wr_idle,

      -- internal interface
      raddr                   => raddr,
      length_bytes            => rlength_bytes,
      rbarhit                 => rbarhit,
      araddr_2lsbs            => araddr_2lsbs,
      last_BE                 => rlast_BE,
      req_active              => rreq_active,
      req_active_ptr          => req_active_ptr,
      read_req_sent           => read_req_sent,
      tag_cpl_status_clr      => tag_cpl_status_clr,
      rdata_bram_rd_en        => rdata_bram_rd_en,
      rdata_bram_addr         => rdata_bram_addr,
      rdata                   => rdata,
      cpl_index               => cpl_index,
      rdata_str_done          => rdata_str_done,
      rdata_str_start         => rdata_str_start,
      first_word_offset       => first_word_offset,
      illegal_burst           => illegal_burst_rd,
      bar_error               => bar_error_rd,
      cpl_timer_timeout_strb  => cpl_timer_timeout_strb,
      unsupported_req         => unsupported_req,
      completer_abort         => completer_abort,
      poisoned_req            => poisoned_req,
      header_ep               => header_ep,
      rd_req_index_err        => rd_req_index_err,
      blk_lnk_up              => blk_lnk_up,
      pcie_bme                => sig_pcie_bme
   );

   -- write data path
   comp_write_data_fifo : xpm_fifo_sync
   generic map (
     FIFO_MEMORY_TYPE         => "block",
     ECC_MODE                 => "no_ecc",
     FIFO_WRITE_DEPTH         => 256,
     WRITE_DATA_WIDTH         => C_S_AXI_DATA_WIDTH,
     WR_DATA_COUNT_WIDTH      => 9,
     PROG_FULL_THRESH         => 10,
     FULL_RESET_VALUE         => 1,
     READ_MODE                => "fwft",
     FIFO_READ_LATENCY        => 0,
     READ_DATA_WIDTH          => C_S_AXI_DATA_WIDTH,
     RD_DATA_COUNT_WIDTH      => 9,
     USE_ADV_FEATURES         => "1F1F",
     PROG_EMPTY_THRESH        => 10,
     DOUT_RESET_VALUE         => "0",
     WAKEUP_TIME              => 0
     )
   port map (
     rst              => reset_inv_wr_fifo,
     wr_clk           => s_axi_aclk,
     wr_en            => wdata_valid1,
     wr_ack           => open,
     din              => wdata1,
     full             => wdata_fifo_full1,
     almost_full      => wdata_fifo_allmost_full1,
     overflow         => open,
     rd_en            => wdata_fifo_rd_en1,
     dout             => wdata_fifo_dout1,
     empty            => wdata_fifo_empty1,
     almost_empty     => open,
     data_valid       => open,
     underflow        => open,
     wr_data_count    => open,
     sleep            => '0',
     injectsbiterr    => '0',
     injectdbiterr    => '0'
     );

   comp_write_data_fifo2 : xpm_fifo_sync
   generic map (
     FIFO_MEMORY_TYPE         => "block",
     ECC_MODE                 => "no_ecc",
     FIFO_WRITE_DEPTH         => 256,
     WRITE_DATA_WIDTH         => C_S_AXI_DATA_WIDTH,
     WR_DATA_COUNT_WIDTH      => 9,
     PROG_FULL_THRESH         => 10,
     FULL_RESET_VALUE         => 1,
     READ_MODE                => "fwft",
     FIFO_READ_LATENCY        => 0,
     READ_DATA_WIDTH          => C_S_AXI_DATA_WIDTH,
     RD_DATA_COUNT_WIDTH      => 9,
     USE_ADV_FEATURES         => "1F1F",
     PROG_EMPTY_THRESH        => 10,
     DOUT_RESET_VALUE         => "0",
     WAKEUP_TIME              => 0
     )
   port map (
     rst              => reset_inv_wr_fifo,
     wr_clk           => s_axi_aclk,
     wr_en            => wdata_valid2,
     wr_ack           => open,
     din              => wdata2,
     full             => wdata_fifo_full2,
     almost_full      => wdata_fifo_allmost_full2,
     overflow         => open,
     rd_en            => wdata_fifo_rd_en2,
     dout             => wdata_fifo_dout2,
     empty            => wdata_fifo_empty2,
     almost_empty     => open,
     data_valid       => open,
     underflow        => open,
     wr_data_count    => open,
     sleep            => '0',
     injectsbiterr    => '0',
     injectdbiterr    => '0'
     );

   -- read data path
   comp_read_data_bram : xpm_memory_tdpram
   generic map (
      MEMORY_SIZE        => (C_S_AXI_DATA_WIDTH * RD_BUFFER_DEPTH),
      MEMORY_PRIMITIVE   => "block",               --string; "auto", "distributed", "block" or "ultra" ;
      CLOCKING_MODE      => "common_clock",
      MEMORY_INIT_FILE   => "none",
      MEMORY_INIT_PARAM  => "",
      USE_MEM_INIT       => 1,
      WAKEUP_TIME        => "disable_sleep",
      MESSAGE_CONTROL    => 0,
      ECC_MODE           => "no_ecc",
      AUTO_SLEEP_TIME    => 0,
      -- Port A module generics
      WRITE_DATA_WIDTH_A => C_S_AXI_DATA_WIDTH,
      READ_DATA_WIDTH_A  => C_S_AXI_DATA_WIDTH,
      BYTE_WRITE_WIDTH_A => 8,
      ADDR_WIDTH_A       => RD_BUFFER_ADDR_SIZE,
      READ_RESET_VALUE_A => "0",
      READ_LATENCY_A     => 1,
      WRITE_MODE_A       => "write_first",
      -- Port B module generics
      WRITE_DATA_WIDTH_B => C_S_AXI_DATA_WIDTH,
      READ_DATA_WIDTH_B  => C_S_AXI_DATA_WIDTH,
      BYTE_WRITE_WIDTH_B => C_S_AXI_DATA_WIDTH,
      ADDR_WIDTH_B       => RD_BUFFER_ADDR_SIZE,
      READ_RESET_VALUE_B => "0",
      READ_LATENCY_B     => 1,
      WRITE_MODE_B       => "write_first"
      )
   port map (
      sleep          => '0',
      -- Port A module ports
      clka           => s_axi_aclk,
      rsta           => '0',   
      ena            => '1',
      regcea         => '1',
      wea            => wea,
      addra          => cpl_buffer_addr,
      dina           => data_stream_out,
      injectsbiterra => '0',
      injectdbiterra => '0',
      douta          => open,
      sbiterra       => open,
      dbiterra       => open,
      -- Port B module ports
      clkb           => s_axi_aclk,
      rstb           => '0',  
      enb            => rdata_bram_rd_en,
      regceb         => '1',
      web            => (OTHERS => '0'),
      addrb          => rdata_bram_addr,
      dinb           => (OTHERS => '0'),
      injectsbiterrb => '0',
      injectdbiterrb => '0',
      doutb          => rdata,
      sbiterrb       => open,
      dbiterrb       => open
      );


-- write streaming interface
   comp_slave_write_req_tlp : entity axi_pcie_v2_9_14.slave_write_req_tlp
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_S_AXI_ADDR_WIDTH      => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH      => C_S_AXI_DATA_WIDTH,
      C_M_AXIS_DATA_WIDTH     => C_M_AXIS_DATA_WIDTH,
      C_AXIBAR_NUM            => C_AXIBAR_NUM,
      C_AXIBAR_0              => C_AXIBAR_0,
      C_AXIBAR_HIGHADDR_0     => C_AXIBAR_HIGHADDR_0,
      C_AXIBAR_1              => C_AXIBAR_1,
      C_AXIBAR_HIGHADDR_1     => C_AXIBAR_HIGHADDR_1,
      C_AXIBAR_2              => C_AXIBAR_2,
      C_AXIBAR_HIGHADDR_2     => C_AXIBAR_HIGHADDR_2,
      C_AXIBAR_3              => C_AXIBAR_3,
      C_AXIBAR_HIGHADDR_3     => C_AXIBAR_HIGHADDR_3,
      C_AXIBAR_4              => C_AXIBAR_4,
      C_AXIBAR_HIGHADDR_4     => C_AXIBAR_HIGHADDR_4,
      C_AXIBAR_5              => C_AXIBAR_5,
      C_AXIBAR_HIGHADDR_5     => C_AXIBAR_HIGHADDR_5,
      C_AXIBAR_AS_0           => C_AXIBAR_AS_0,
      C_AXIBAR_AS_1           => C_AXIBAR_AS_1,
      C_AXIBAR_AS_2           => C_AXIBAR_AS_2,
      C_AXIBAR_AS_3           => C_AXIBAR_AS_3,
      C_AXIBAR_AS_4           => C_AXIBAR_AS_4,
      C_AXIBAR_AS_5           => C_AXIBAR_AS_5,
      C_AXIBAR_CHK_SLV_ERR    => C_AXIBAR_CHK_SLV_ERR
   )
   port map(

      -- AXI Global
      aclk                    => s_axi_aclk,
      reset                   => reset,

      -- internal interface
      maxpayloadsize          => maxpayloadsize,
      waddr                   => waddr,
      length_bytes            => wlength_bytes,
      wbarhit                 => wbarhit,
      wdata                   => wdata_fifo_dout,
      first_BE                => wfirst_BE,
      first_BE_valid          => wfirst_BE_valid,
      last_BE                 => wlast_BE,
      last_BE_valid           => wlast_BE_valid,
      first_word_offset       => wfirst_word_offset,
      wdata_fifo_rd_en        => wdata_fifo_rd_en,
      wdata_fifo_empty        => wdata_fifo_empty,
      reqID                   => reqID,
      wdata_str_done          => wdata_str_done,
      wdata_str_start         => wdata_str_start,
      illegal_burst_trns      => illegal_burst_trns_wr,
      bar_error_trns          => bar_error_trns_wr,
      block_trns_lnkdwn       => block_trns_lnkdwn,
      blk_lnk_up              => blk_lnk_up,
      pcie_bme                => sig_pcie_bme,
      tlp_str_start           => sig_tlp_str_start,

      -- AXI2PCIE translation vectors
      axibar2pciebar0         => axibar2pciebar0,
      axibar2pciebar1         => axibar2pciebar1,
      axibar2pciebar2         => axibar2pciebar2,
      axibar2pciebar3         => axibar2pciebar3,
      axibar2pciebar4         => axibar2pciebar4,
      axibar2pciebar5         => axibar2pciebar5,

      -- AXI Streaming interface
      m_axis_rw_tvalid        => sig_m_axis_rw_tvalid,
      m_axis_rw_tready        => m_axis_rw_tready,
      m_axis_rw_tdata         => m_axis_rw_tdata,
      m_axis_rw_tstrb         => m_axis_rw_tstrb,
      m_axis_rw_tlast         => m_axis_rw_tlast
   );


-- read request streaming interface
   comp_slave_read_req_tlp : entity axi_pcie_v2_9_14.slave_read_req_tlp
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_S_AXI_ID_WIDTH        => C_S_AXI_ID_WIDTH,
      C_S_AXI_ADDR_WIDTH      => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH      => C_S_AXI_DATA_WIDTH,
      C_M_AXIS_DATA_WIDTH     => C_M_AXIS_DATA_WIDTH,
      C_AXIBAR_NUM            => C_AXIBAR_NUM,
      C_AXIBAR_0              => C_AXIBAR_0,
      C_AXIBAR_HIGHADDR_0     => C_AXIBAR_HIGHADDR_0,
      C_AXIBAR_1              => C_AXIBAR_1,
      C_AXIBAR_HIGHADDR_1     => C_AXIBAR_HIGHADDR_1,
      C_AXIBAR_2              => C_AXIBAR_2,
      C_AXIBAR_HIGHADDR_2     => C_AXIBAR_HIGHADDR_2,
      C_AXIBAR_3              => C_AXIBAR_3,
      C_AXIBAR_HIGHADDR_3     => C_AXIBAR_HIGHADDR_3,
      C_AXIBAR_4              => C_AXIBAR_4,
      C_AXIBAR_HIGHADDR_4     => C_AXIBAR_HIGHADDR_4,
      C_AXIBAR_5              => C_AXIBAR_5,
      C_AXIBAR_HIGHADDR_5     => C_AXIBAR_HIGHADDR_5,
      C_AXIBAR_AS_0           => C_AXIBAR_AS_0,
      C_AXIBAR_AS_1           => C_AXIBAR_AS_1,
      C_AXIBAR_AS_2           => C_AXIBAR_AS_2,
      C_AXIBAR_AS_3           => C_AXIBAR_AS_3,
      C_AXIBAR_AS_4           => C_AXIBAR_AS_4,
      C_AXIBAR_AS_5           => C_AXIBAR_AS_5,
      C_EP_LINK_PARTNER_RCB   => C_EP_LINK_PARTNER_RCB
   )
   port map(

      -- AXI Global
      aclk                    => s_axi_aclk,
      reset                   => reset,

      -- internal interface
      maxreadreqsize          => maxreadreqsize,
      raddr                   => raddr,
      length_bytes            => rlength_bytes,
      rbarhit                 => rbarhit,
      araddr_2lsbs            => araddr_2lsbs,
      last_BE                 => rlast_BE,
      reqID                   => reqID,
      req_active              => rreq_active,
      read_req_sent           => read_req_sent,
      tag_sent                => tag_sent,
      length_sent             => length_sent,
      illegal_burst           => illegal_burst_rd,
      illegal_burst_trns      => illegal_burst_trns_rd,
      bar_error               => bar_error_rd,
      bar_error_trns          => bar_error_trns_rd,
      total_length_out        => total_length_out,
      pcie_bme                => sig_pcie_bme,
      blk_lnk_up              => blk_lnk_up,
      tag_pending_for_cpl     => tag_pending_for_cpl,

      -- AXI2PCIE translation vectors
      axibar2pciebar0         => axibar2pciebar0,
      axibar2pciebar1         => axibar2pciebar1,
      axibar2pciebar2         => axibar2pciebar2,
      axibar2pciebar3         => axibar2pciebar3,
      axibar2pciebar4         => axibar2pciebar4,
      axibar2pciebar5         => axibar2pciebar5,

      -- AXI Streaming interface
      m_axis_rr_tvalid        => sig_m_axis_rr_tvalid,
      m_axis_rr_tready        => m_axis_rr_tready,
      m_axis_rr_tdata         => m_axis_rr_tdata,
      m_axis_rr_tstrb         => m_axis_rr_tstrb,
      m_axis_rr_tlast         => sig_m_axis_rr_tlast,
      config_gen_req          => config_gen_req
   );


-- read completions streaming interface
   comp_slave_read_cpl_tlp : entity axi_pcie_v2_9_14.slave_read_cpl_tlp
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_AXIREAD_NUM           => C_AXIREAD_NUM,
      C_RD_BUFFER_ADDR_SIZE   => RD_BUFFER_ADDR_SIZE,
      C_M_AXIS_DATA_WIDTH     => C_M_AXIS_DATA_WIDTH
   )
   port map(
      -- AXI Global
      aclk                    => s_axi_aclk,
      reset                   => reset,

      -- internal interface
      maxreadreqsize          => maxreadreqsize,--: in  std_logic_vector(2 downto 0);
      m_axis_rr_tlast         => sig_m_axis_rr_tlast,
      m_axis_rr_tready        => m_axis_rr_tready,
      read_req_sent           => read_req_sent,
      tag_sent                => tag_sent,--: in  std_logic_vector(7 downto 0);
      length_sent             => length_sent,--: in  std_logic_vector(9 downto 0);
      rreq_active             => rreq_active,--: in  std_logic;
      req_active_ptr          => req_active_ptr,--: in  integer range 0 to 7;
      data_stream_out         => data_stream_out,--: out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      read_data_bram_we       => wea,--: out std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
      cpl_buffer_addr         => cpl_buffer_addr,--: out std_logic_vector(10 downto 0);
      cpl_data_str_done       => cpl_data_str_done,--: out std_logic;
      tag_in_cpl              => tag_in_cpl,--: out std_logic_vector(7 downto 0);
      tag_cpl_status_clr      => tag_cpl_status_clr,
      cpl_index               => cpl_index,
      rdata_str_done          => rdata_str_done,
      rdata_str_start         => rdata_str_start,
      first_word_offset       => first_word_offset,
      unsupported_req         => unsupported_req,
      completer_abort         => completer_abort,
      poisoned_req            => poisoned_req,
      unexpected_cpl          => unexpected_cpl,
      cpl_timer_timeout_strb  => cpl_timer_timeout_strb,
      rd_req_index_err        => rd_req_index_err,
      blk_lnk_up              => blk_lnk_up,
      header_ep               => header_ep,
      reqID                   => reqID,
      illegal_burst_trns      => illegal_burst_trns_rd,
      bar_error_trns          => bar_error_trns_rd,
      total_length_out        => total_length_out,
      tag_pending_for_cpl     => tag_pending_for_cpl,
      tag_len_active_valid_o  => tag_len_active_valid,

      -- AXI Streaming interface
      s_axis_rc_tdata         => s_axis_rc_tdata,--: in  std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      s_axis_rc_tstrb         => s_axis_rc_tstrb,--: in  std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      s_axis_rc_tlast         => s_axis_rc_tlast,--: in  std_logic;
      s_axis_rc_tvalid        => s_axis_rc_tvalid,--: in  std_logic;
      s_axis_rc_tready        => s_axis_rc_tready--: out std_logic
   );



gen_axi_upsizer : if C_S_AXI_SUPPORTS_NARROW_BURST = 1 generate



-- axi_upsizer implemented
comp_axi_upsizer : axi_pcie_v2_9_14_axi_upsizer
    generic map(
        C_FAMILY                    => "rtl",            --: string  := "none";
        C_AXI_ID_WIDTH              => C_S_AXI_ID_WIDTH,    --: integer := 4;
        C_AXI_ADDR_WIDTH            => C_S_AXI_ADDR_WIDTH,  --: integer := 32;
        C_S_AXI_DATA_WIDTH          => C_S_AXI_DATA_WIDTH,  --: integer := 32;
        C_M_AXI_DATA_WIDTH          => C_S_AXI_DATA_WIDTH,  --: integer := 64;
        C_AXI_SUPPORTS_WRITE        => 1,                   --: integer := 1;
        C_AXI_SUPPORTS_READ         => 1,                   --: integer := 1;
        C_S_AXI_R_REGISTER          => 0,                -- CR # 649227
        C_M_AXI_R_REGISTER          => 0,                -- CR # 649227
        C_PACKING_LEVEL             => 2,                   --: integer := 1;
        C_SUPPORT_BURSTS            => 1,                   --: integer := 1;
        C_SINGLE_THREAD             => 0                    --: integer := 1
    )
    port map(
   -- Globals
        ARESETN                     => reset,              --:in  std_logic;
        ACLK                        => s_axi_aclk,         --:in  std_logic;
   -- Slave Interface Write Address Ports
        S_AXI_AWID                  => s_axi_awid,         --:in  std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        S_AXI_AWADDR                => s_axi_awaddr,       --:in  std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
        S_AXI_AWLEN                 => s_axi_awlen,        --:in  std_logic_vector(7 downto 0);
        S_AXI_AWSIZE                => s_axi_awsize,       --:in  std_logic_vector(2 downto 0);
        S_AXI_AWBURST               => s_axi_awburst,      --:in  std_logic_vector(1 downto 0);
        S_AXI_AWLOCK                => "00",               --:in  std_logic_vector(1 downto 0);
        S_AXI_AWCACHE               => "0000",             --:in  std_logic_vector(3 downto 0);
        S_AXI_AWPROT                => "000",              --:in  std_logic_vector(2 downto 0);
        S_AXI_AWREGION              => s_axi_awregion,     --:in  std_logic_vector(3 downto 0);
        S_AXI_AWQOS                 => "0000",             --:in  std_logic_vector(3 downto 0);
        S_AXI_AWUSER                => "0",                --:in  std_logic_vector(C_AXI_AWUSER_WIDTH-1 downto 0);
        S_AXI_AWVALID               => s_axi_awvalid,      --:in  std_logic;
        S_AXI_AWREADY               => s_axi_awready,      --:out std_logic;
   -- Slave Interface Write Data Ports
        S_AXI_WDATA                 => s_axi_wdata,        --:in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
        S_AXI_WSTRB                 => s_axi_wstrb,        --:in  std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
        S_AXI_WLAST                 => s_axi_wlast,        --:in  std_logic;
        S_AXI_WUSER                 => "0",                --:in  std_logic_vector(C_AXI_WUSER_WIDTH-1 downto 0);
        S_AXI_WVALID                => s_axi_wvalid,       --:in  std_logic;
        S_AXI_WREADY                => s_axi_wready,       --:out std_logic;
   -- Slave Interface Write Response Ports
        S_AXI_BID                   => s_axi_bid,          --:out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        S_AXI_BRESP                 => s_axi_bresp,        --:out std_logic_vector(1 downto 0);
        S_AXI_BVALID                => s_axi_bvalid,       --:out std_logic;
        S_AXI_BREADY                => s_axi_bready,       --:in  std_logic;
   -- Slave Interface Read Address Ports
        S_AXI_ARID                  => s_axi_arid,         --:in  std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        S_AXI_ARADDR                => s_axi_araddr,       --:in  std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
        S_AXI_ARLEN                 => s_axi_arlen,        --:in  std_logic_vector(7 downto 0);
        S_AXI_ARSIZE                => s_axi_arsize,       --:in  std_logic_vector(2 downto 0);
        S_AXI_ARBURST               => s_axi_arburst,      --:in  std_logic_vector(1 downto 0);
        S_AXI_ARLOCK                => "00",               --:in  std_logic_vector(1 downto 0);
        S_AXI_ARCACHE               => "0000",             --:in  std_logic_vector(3 downto 0);
        S_AXI_ARPROT                => "000",              --:in  std_logic_vector(2 downto 0);
        S_AXI_ARREGION              => s_axi_arregion,     --:in  std_logic_vector(3 downto 0);
        S_AXI_ARQOS                 => "0000",             --:in  std_logic_vector(3 downto 0);
        S_AXI_ARUSER                => "0",                --:in  std_logic_vector(C_AXI_ARUSER_WIDTH-1 downto 0);
        S_AXI_ARVALID               => s_axi_arvalid,      --:in  std_logic;
        S_AXI_ARREADY               => sig_s_axi_arready,  --:out std_logic;
   -- Slave Interface Read Data Ports
        S_AXI_RID                   => s_axi_rid,          --:out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        S_AXI_RDATA                 => s_axi_rdata,        --:out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
        S_AXI_RRESP                 => s_axi_rresp,        --:out std_logic_vector(1 downto 0);
        S_AXI_RLAST                 => s_axi_rlast,        --:out std_logic;
        S_AXI_RVALID                => s_axi_rvalid,       --:out std_logic;
        S_AXI_RREADY                => s_axi_rready,       --:in  std_logic;
   -- Master Interface Write Address Port
        M_AXI_AWID                  => sig_m_axi_awid,     --:out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        M_AXI_AWADDR                => sig_m_axi_awaddr,   --:out std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
        M_AXI_AWLEN                 => sig_m_axi_awlen,    --:out std_logic_vector(7 downto 0);
        M_AXI_AWSIZE                => sig_m_axi_awsize,   --:out std_logic_vector(2 downto 0);
        M_AXI_AWBURST               => sig_m_axi_awburst,  --:out std_logic_vector(1 downto 0);
        M_AXI_AWREGION              => sig_m_axi_awregion, --:out std_logic_vector(3 downto 0);
        M_AXI_AWVALID               => sig_m_axi_awvalid,  --:out std_logic;
        M_AXI_AWREADY               => sig_m_axi_awready,  --:in  std_logic;
   -- Master Interface Write Data Ports
        M_AXI_WDATA                 => sig_m_axi_wdata,    --:out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
        M_AXI_WSTRB                 => sig_m_axi_wstrb,    --:out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0);
        M_AXI_WLAST                 => sig_m_axi_wlast,    --:out std_logic;
        M_AXI_WVALID                => sig_m_axi_wvalid,   --:out std_logic;
        M_AXI_WREADY                => sig_m_axi_wready,   --:in  std_logic;
   -- Master Interface Write Response Ports
        M_AXI_BID                   => sig_m_axi_bid,      --:in  std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        M_AXI_BRESP                 => sig_m_axi_bresp,    --:in  std_logic_vector(1 downto 0);
        M_AXI_BUSER                 => "0",                --:in  std_logic_vector(C_AXI_BUSER_WIDTH-1 downto 0);
        M_AXI_BVALID                => sig_m_axi_bvalid,   --:in  std_logic;
        M_AXI_BREADY                => sig_m_axi_bready,   --:out std_logic;
   -- Master Interface Read Address Port
        M_AXI_ARID                  => sig_m_axi_arid,     --:out std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        M_AXI_ARADDR                => sig_m_axi_araddr,   --:out std_logic_vector(C_AXI_ADDR_WIDTH-1 downto 0);
        M_AXI_ARLEN                 => sig_m_axi_arlen,    --:out std_logic_vector(7 downto 0);
        M_AXI_ARSIZE                => sig_m_axi_arsize,   --:out std_logic_vector(2 downto 0);
        M_AXI_ARBURST               => sig_m_axi_arburst,  --:out std_logic_vector(1 downto 0);
        M_AXI_ARREGION              => sig_m_axi_arregion, --:out std_logic_vector(3 downto 0);
        M_AXI_ARVALID               => sig_m_axi_arvalid,  --:out std_logic;
        M_AXI_ARREADY               => sig_m_axi_arready,  --:in  std_logic;
   -- Master Interface Read Data Ports
        M_AXI_RID                   => sig_m_axi_rid,      --:in  std_logic_vector(C_AXI_ID_WIDTH-1 downto 0);
        M_AXI_RDATA                 => sig_m_axi_rdata,    --:in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
        M_AXI_RRESP                 => sig_m_axi_rresp,    --:in  std_logic_vector(1 downto 0);
        M_AXI_RLAST                 => sig_m_axi_rlast,    --:in  std_logic;
        M_AXI_RUSER                 => "0",                --:in  std_logic_vector(C_AXI_RUSER_WIDTH-1 downto 0);
        M_AXI_RVALID                => sig_m_axi_rvalid,   --:in  std_logic;
        M_AXI_RREADY                => sig_m_axi_rready    --:out std_logic
   );

   s_axi_arready  <= sig_s_axi_arready;
   pu_axi_arsize_len_sync : process (s_axi_aclk)
   begin
      if (rising_edge(s_axi_aclk)) then
         if reset = '0' then
            pu_axi_arlen_d  <= (others => '0');
            pu_axi_arsize_d <= (others => '0');
         elsif s_axi_arvalid = '1' and sig_s_axi_arready = '1' then
            pu_axi_arlen_d  <= s_axi_arlen;
            pu_axi_arsize_d <= s_axi_arsize;
         end if;
      end if;
   end process;
end generate;

gen_no_axi_upsizer : if C_S_AXI_SUPPORTS_NARROW_BURST = 0 generate

-- no axi_upsizer implemented

   -- Slave Interface Write Address Ports
   sig_m_axi_awid                  <= s_axi_awid;
   sig_m_axi_awaddr                <= s_axi_awaddr;
   sig_m_axi_awlen                 <= s_axi_awlen;
   sig_m_axi_awsize                <= s_axi_awsize;
   sig_m_axi_awburst               <= s_axi_awburst;
   sig_m_axi_awregion              <= s_axi_awregion;
   sig_m_axi_awvalid               <= s_axi_awvalid;
   s_axi_awready                   <= sig_m_axi_awready;
   -- Slave Interface Write Data Ports
   sig_m_axi_wdata                 <= s_axi_wdata;
   sig_m_axi_wstrb                 <= s_axi_wstrb;
   sig_m_axi_wlast                 <= s_axi_wlast;
   sig_m_axi_wvalid                <= s_axi_wvalid;
   s_axi_wready                    <= sig_m_axi_wready;
   -- Slave Interface Write Response Ports
   s_axi_bid                       <= sig_m_axi_bid;
   s_axi_bresp                     <= sig_m_axi_bresp;
   s_axi_bvalid                    <= sig_m_axi_bvalid;
   sig_m_axi_bready                <= s_axi_bready;
   -- Slave Interface Read Address Ports
   sig_m_axi_arid                  <= s_axi_arid;
   sig_m_axi_araddr                <= s_axi_araddr;
   sig_m_axi_arlen                 <= s_axi_arlen;
   sig_m_axi_arsize                <= s_axi_arsize;
   sig_m_axi_arburst               <= s_axi_arburst;
   sig_m_axi_arregion              <= s_axi_arregion;
   sig_m_axi_arvalid               <= s_axi_arvalid;
   s_axi_arready                   <= sig_m_axi_arready;
   -- Slave Interface Read Data Ports
   s_axi_rid                       <= sig_m_axi_rid;
   s_axi_rdata                     <= sig_m_axi_rdata;
   s_axi_rresp                     <= sig_m_axi_rresp;
   s_axi_rlast                     <= sig_m_axi_rlast;
   s_axi_rvalid                    <= sig_m_axi_rvalid;
   sig_m_axi_rready                <= s_axi_rready;
   -- pre-upsizer signals
   pu_axi_arlen_d                  <= s_axi_arlen;
   pu_axi_arsize_d                 <= s_axi_arsize;

end generate;


end architecture;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_pcie_mm_s.vhd
--
-- Description:     Ensure the Bar hit for RP & EP configuration 
--        is incorporated between this bridge core and 
--        enhanced PCIe core.
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--              axi_pcie_mm_s.vhd
--
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;

library axi_pcie_v2_9_14;

--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------



entity axi_pcie_mm_s is
   generic(
      --Family Generics
      C_FAMILY                      : string; --  :="virtex7";
      C_S_AXI_ID_WIDTH              : integer; -- := 4;
      --C_M_AXI_THREAD_ID_WIDTH       : integer; -- := 4;
      C_S_AXI_ADDR_WIDTH            : integer; -- := 32;
      C_S_AXI_DATA_WIDTH            : integer; -- := 32;
      C_M_AXI_ADDR_WIDTH            : integer; -- := 32;
      C_M_AXI_DATA_WIDTH            : integer; -- := 32;
      C_S_AXIS_DATA_WIDTH           : integer; -- := 32;
      C_M_AXIS_DATA_WIDTH           : integer; -- := 32;
      C_COMP_TIMEOUT                : integer; -- := 0;
      C_USER_CLK_FREQ               : integer; -- := 1;
      C_USER_CLK2_DIV2              : string;  -- := "FALSE";
      C_INCLUDE_RC                  : integer; -- := 0;
      C_S_AXI_SUPPORTS_NARROW_BURST : integer; -- := 1;
      C_EP_LINK_PARTNER_RCB         : integer := 0;
      C_INCLUDE_BAROFFSET_REG       : integer; -- := 1;
      C_AXIREAD_NUM                 : integer := 8;    -- CR # 646225
      C_AXIBAR_NUM                  : integer; -- := 6;
      C_AXIBAR2PCIEBAR_0            : std_logic_vector; --:=x"00000000";
      C_AXIBAR2PCIEBAR_1            : std_logic_vector; --:=x"00000000";
      C_AXIBAR2PCIEBAR_2            : std_logic_vector; --:=x"00000000";
      C_AXIBAR2PCIEBAR_3            : std_logic_vector; --:=x"00000000";
      C_AXIBAR2PCIEBAR_4            : std_logic_vector; --:=x"00000000";
      C_AXIBAR2PCIEBAR_5            : std_logic_vector; --:=x"00000000";
      C_AXIBAR_AS_0                 : integer; -- := 0;
      C_AXIBAR_AS_1                 : integer; -- := 0;
      C_AXIBAR_AS_2                 : integer; -- := 0;
      C_AXIBAR_AS_3                 : integer; -- := 0;
      C_AXIBAR_AS_4                 : integer; -- := 0;
      C_AXIBAR_AS_5                 : integer; -- := 0;
      C_AXIBAR_0                    : std_logic_vector; -- := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0           : std_logic_vector; -- := x"0000_0000";
      C_AXIBAR_1                    : std_logic_vector; -- := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1           : std_logic_vector; -- := x"0000_0000";
      C_AXIBAR_2                    : std_logic_vector; -- := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2           : std_logic_vector; -- := x"0000_0000";
      C_AXIBAR_3                    : std_logic_vector; -- := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3           : std_logic_vector; -- := x"0000_0000";
      C_AXIBAR_4                    : std_logic_vector; -- := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4           : std_logic_vector; -- := x"0000_0000";
      C_AXIBAR_5                    : std_logic_vector; -- := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5           : std_logic_vector; -- := x"0000_0000";
      C_PCIEBAR_NUM                 : integer; -- := 3;
      C_PCIEBAR_AS                  : integer; -- := 1;
      C_PCIEBAR_LEN_0               : integer; -- := 16;
      C_PCIEBAR2AXIBAR_0            : std_logic_vector; --:=x"00000000";
      C_PCIEBAR2AXIBAR_0_SEC        : integer; -- := 0;
      C_PCIEBAR_LEN_1               : integer; -- := 16;
      C_PCIEBAR2AXIBAR_1            : std_logic_vector; --:=x"00000000";
      C_PCIEBAR2AXIBAR_1_SEC        : integer; -- := 0;
      C_PCIEBAR_LEN_2               : integer; -- := 16;
      C_PCIEBAR2AXIBAR_2            : std_logic_vector; --:=x"00000000";
      C_PCIEBAR2AXIBAR_2_SEC        : integer; -- := 0;
      C_S_AXIS_USER_WIDTH           : integer; -- := 12;
      C_TRN_NP_FC                   : string;   -- := "FALSE";
      C_AXIBAR_CHK_SLV_ERR          : string   -- := "FALSE"
      --C_M_AXI_AWUSER_WIDTH    : integer;
      --C_M_AXI_WUSER_WIDTH     : integer
      --C_NUM_USER_INTR         : integer := 6
   );
   port(

      -- AXI Global
      axi_aclk                : in  std_logic;
      reset                   : in  std_logic;

      -- AXI Slave Write Address Channel
      s_axi_awid              : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_awaddr            : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_awregion          : in  std_logic_vector(3 downto 0);
      s_axi_awlen             : in  std_logic_vector(7 downto 0);
      s_axi_awsize            : in  std_logic_vector(2 downto 0);
      s_axi_awburst           : in  std_logic_vector(1 downto 0);
      s_axi_awvalid           : in  std_logic;
      s_axi_awready           : out std_logic;

      -- AXI Slave Write Data Channel
      s_axi_wdata             : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_wstrb             : in  std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
      s_axi_wlast             : in  std_logic;
      s_axi_wvalid            : in  std_logic;
      s_axi_wready            : out std_logic;

      -- AXI Slave Write Response Channel
      s_axi_bid               : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_bresp             : out std_logic_vector(1 downto 0);
      s_axi_bvalid            : out std_logic;
      s_axi_bready            : in  std_logic;

      -- AXI Slave Read Address Channel
      s_axi_arid              : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_araddr            : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_arregion          : in  std_logic_vector(3 downto 0);
      s_axi_arlen             : in  std_logic_vector(7 downto 0);
      s_axi_arsize            : in  std_logic_vector(2 downto 0);
      s_axi_arburst           : in  std_logic_vector(1 downto 0);
      s_axi_arvalid           : in  std_logic;
      s_axi_arready           : out std_logic;

      -- AXI Slave Read Data Channel
      s_axi_rid               : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_rdata             : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_rresp             : out std_logic_vector(1 downto 0);
      s_axi_rlast             : out std_logic;
      s_axi_rvalid            : out std_logic;
      s_axi_rready            : in  std_logic;

      -- AXIS Write Requester Channel
      m_axis_rw_tdata         : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_rw_tstrb         : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_rw_tlast         : out std_logic;
      m_axis_rw_tvalid        : out std_logic;
      m_axis_rw_tready        : in  std_logic;

      -- AXIS Read Requester Channel
      m_axis_rr_tid           : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      m_axis_rr_tdata         : out std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_rr_tstrb         : out std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_rr_tlast         : out std_logic;
      m_axis_rr_tvalid        : out std_logic;
      m_axis_rr_tready        : in  std_logic;

      -- AXIS Completion Requester Channel
      s_axis_rc_tdata         : in  std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
      s_axis_rc_tstrb         : in  std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
      s_axis_rc_tlast         : in  std_logic;
      s_axis_rc_tvalid        : in  std_logic;
      s_axis_rc_tready        : out std_logic;

      -- AXI Master Write Address Channel
      m_axi_awaddr            : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
      m_axi_awlen             : out std_logic_vector(7 downto 0);
      m_axi_awsize            : out std_logic_vector(2 downto 0);
      m_axi_awburst           : out std_logic_vector(1 downto 0);
      m_axi_awprot            : out std_logic_vector(2 downto 0);
      m_axi_awvalid           : out std_logic;
      m_axi_awready           : in  std_logic;
      --m_axi_awid              : out std_logic_vector(C_M_AXI_THREAD_ID_WIDTH-1 downto 0);
      m_axi_awlock            : out std_logic;
      m_axi_awcache           : out std_logic_vector(3 downto 0);

      -- AXI Master Write Data Channel
      m_axi_wdata             : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
      m_axi_wstrb             : out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0);
      m_axi_wlast             : out std_logic;
      m_axi_wvalid            : out std_logic;
      m_axi_wready            : in  std_logic;

      -- AXI Master Write Response Channel
      m_axi_bresp             : in  std_logic_vector(1 downto 0);
      m_axi_bvalid            : in  std_logic;
      m_axi_bready            : out std_logic;

      -- AXI Master Read Address Channel
      --m_axi_arid              : out std_logic_vector(C_M_AXI_THREAD_ID_WIDTH-1 downto 0);
      m_axi_araddr            : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
      m_axi_arlen             : out std_logic_vector(7 downto 0);
      m_axi_arsize            : out std_logic_vector(2 downto 0);
      m_axi_arburst           : out std_logic_vector(1 downto 0);
      m_axi_arprot            : out std_logic_vector(2 downto 0);
      m_axi_arvalid           : out std_logic;
      m_axi_arready           : in  std_logic;
      m_axi_arlock            : out std_logic;
      m_axi_arcache           : out std_logic_vector(3 downto 0);
      --m_axi_aruser            : out std_logic_vector(C_M_AXI_AWUSER_WIDTH-1 downto 0);

      -- AXI Master Read Data Channel
      m_axi_rdata             : in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
      m_axi_rresp             : in  std_logic_vector(1 downto 0);
      m_axi_rlast             : in  std_logic;
      m_axi_rvalid            : in  std_logic;
      m_axi_rready            : out std_logic;
      --m_axi_ruser             : out std_logic_vector(C_M_AXI_WUSER_WIDTH-1 downto 0);

      -- AXIS Write Completer Channel
      s_axis_cw_tdata         : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
      s_axis_cw_tstrb         : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
      s_axis_cw_tlast         : in  std_logic;
      s_axis_cw_tvalid        : in  std_logic;
      s_axis_cw_tready        : out std_logic;
      s_axis_cw_tuser         : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0);
      
      -- AXIS Read Completer Channel
      s_axis_cr_tdata         : in  std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
      s_axis_cr_tstrb         : in  std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
      s_axis_cr_tlast         : in  std_logic;
      s_axis_cr_tvalid        : in  std_logic;
      s_axis_cr_tready        : out std_logic;
      s_axis_cr_tuser         : in  std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0);

      -- AXIS Completion Completer Channel
      m_axis_cc_tdata         : out std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
      m_axis_cc_tstrb         : out std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
      m_axis_cc_tlast         : out std_logic;
      m_axis_cc_tvalid        : out std_logic;
      m_axis_cc_tready        : in  std_logic;
      m_axis_cc_tuser         : out std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0);

      -- AXI-Lite Slave IPIC
      IP2Bus_Data             : out std_logic_vector(31 downto 0);
      IP2Bus_WrAck            : out std_logic;
      IP2Bus_RdAck            : out std_logic;
      IP2Bus_Error            : out std_logic;
      Bus2IP_Addr             : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      Bus2IP_Data             : in  std_logic_vector(31 downto 0);
      Bus2IP_RNW              : in  std_logic;
      Bus2IP_BE               : in  std_logic_vector(32/8-1 downto 0);
      Bus2IP_CS               : in  std_logic;

      -- AXI-S Block Interface
      blk_lnk_up              : in  std_logic;
      blk_bus_number          : in  std_logic_vector(7 downto 0);
      blk_device_number       : in  std_logic_vector(4 downto 0);
      blk_function_number     : in  std_logic_vector(2 downto 0);
      blk_command             : in  std_logic_vector(15 downto 0);
      blk_dcontrol            : in  std_logic_vector(15 downto 0);
      blk_lstatus             : in  std_logic_vector(15 downto 0);
      np_cpl_pending          : out std_logic;
      RP_bridge_en            : in  std_logic;

      --Interrupt Strobes
      SUR_int                 : out std_logic;
      SUC_int                 : out std_logic;
      SCT_int                 : out std_logic;
      SEP_int                 : out std_logic;
      SCA_int                 : out std_logic;
      SIB_int                 : out std_logic;
      MDE_int                 : out std_logic; -- Master DECERR interrupt
      MSE_int                 : out std_logic; -- Master SLVERR interrupt
      MEP_int                 : out std_logic; -- Slave Error Poison interrupt
      --MLE_int                 : out std_logic; -- Link Down interrupt
      --MEC_int                 : out std_logic  -- ECRC Error interrupt
      -- signals used to keep track NP buffer availability
      rdndreqpipeline         : out std_logic_vector(2 downto 0);
      rdreqpipeline           : out std_logic_vector(2 downto 0);
      np_pkt_complete         : out std_logic_vector(1 downto 0);
      config_gen_req          : in  std_logic
   );

end axi_pcie_mm_s;

architecture structure of axi_pcie_mm_s is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";

   signal axibar2pciebar0     : std_logic_vector(63 downto 0);
   signal axibar2pciebar1     : std_logic_vector(63 downto 0);
   signal axibar2pciebar2     : std_logic_vector(63 downto 0);
   signal axibar2pciebar3     : std_logic_vector(63 downto 0);
   signal axibar2pciebar4     : std_logic_vector(63 downto 0);
   signal axibar2pciebar5     : std_logic_vector(63 downto 0);
   
   signal slwrreqpendsig              : std_logic_vector(1 downto 0);
   signal slwrreqcompsig              : std_logic_vector(1 downto 0);
   signal sig_slv_write_idle          : std_logic;
   signal sig_s_axi_awvalid           : std_logic;
   signal sig_master_wr_idle          : std_logic;
   signal wrreqpendsig, wrreqcompsig  : std_logic_vector(2 downto 0);
   
begin

   comp_register_block : entity axi_pcie_v2_9_14.register_block
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      C_S_AXI_ADDR_WIDTH      => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH      => C_S_AXI_DATA_WIDTH,
      C_AXIBAR_NUM            => C_AXIBAR_NUM,
      C_INCLUDE_BAROFFSET_REG => C_INCLUDE_BAROFFSET_REG,
      C_AXIBAR2PCIEBAR_0      => C_AXIBAR2PCIEBAR_0,
      C_AXIBAR2PCIEBAR_1      => C_AXIBAR2PCIEBAR_1,
      C_AXIBAR2PCIEBAR_2      => C_AXIBAR2PCIEBAR_2,
      C_AXIBAR2PCIEBAR_3      => C_AXIBAR2PCIEBAR_3,
      C_AXIBAR2PCIEBAR_4      => C_AXIBAR2PCIEBAR_4,
      C_AXIBAR2PCIEBAR_5      => C_AXIBAR2PCIEBAR_5,
      C_AXIBAR_AS_0           => C_AXIBAR_AS_0,
      C_AXIBAR_AS_1           => C_AXIBAR_AS_1,
      C_AXIBAR_AS_2           => C_AXIBAR_AS_2,
      C_AXIBAR_AS_3           => C_AXIBAR_AS_3,
      C_AXIBAR_AS_4           => C_AXIBAR_AS_4,
      C_AXIBAR_AS_5           => C_AXIBAR_AS_5
   )
   port map(
      -- AXI Global
      s_axi_aclk              => axi_aclk,
      reset                   => reset,

      -- AXI-Lite Slave IPIC
      IP2Bus_Data             => IP2Bus_Data,
      IP2Bus_WrAck            => IP2Bus_WrAck,
      IP2Bus_RdAck            => IP2Bus_RdAck,
      IP2Bus_Error            => IP2Bus_Error,
      Bus2IP_Addr             => Bus2IP_Addr,
      Bus2IP_Data             => Bus2IP_Data,
      Bus2IP_RNW              => Bus2IP_RNW,
      Bus2IP_BE               => Bus2IP_BE,
      Bus2IP_CS               => Bus2IP_CS,
      axibar2pciebar0         => axibar2pciebar0,
      axibar2pciebar1         => axibar2pciebar1,
      axibar2pciebar2         => axibar2pciebar2,
      axibar2pciebar3         => axibar2pciebar3,
      axibar2pciebar4         => axibar2pciebar4,
      axibar2pciebar5         => axibar2pciebar5
   );

comp_AXI_MM_S_MasterBridge: entity axi_pcie_v2_9_14.AXI_MM_S_MasterBridge
   generic map(
      --Family Generics
      C_FAMILY                => C_FAMILY,
      --C_M_AXI_THREAD_ID_WIDTH => C_M_AXI_THREAD_ID_WIDTH,
      C_M_AXI_ADDR_WIDTH      => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH      => C_M_AXI_DATA_WIDTH,
      C_S_AXIS_DATA_WIDTH     => C_S_AXIS_DATA_WIDTH,
      C_PCIEBAR_NUM           => C_PCIEBAR_NUM,
      C_PCIEBAR_AS            => C_PCIEBAR_AS,
      C_PCIEBAR_LEN_0         => C_PCIEBAR_LEN_0,
      C_PCIEBAR2AXIBAR_0      => C_PCIEBAR2AXIBAR_0,
      C_PCIEBAR2AXIBAR_0_SEC  => C_PCIEBAR2AXIBAR_0_SEC,
      C_PCIEBAR_LEN_1         => C_PCIEBAR_LEN_1,
      C_PCIEBAR2AXIBAR_1      => C_PCIEBAR2AXIBAR_1,
      C_PCIEBAR2AXIBAR_1_SEC  => C_PCIEBAR2AXIBAR_1_SEC,
      C_PCIEBAR_LEN_2         => C_PCIEBAR_LEN_2,
      C_PCIEBAR2AXIBAR_2      => C_PCIEBAR2AXIBAR_2,
      C_PCIEBAR2AXIBAR_2_SEC  => C_PCIEBAR2AXIBAR_2_SEC,
      C_S_AXIS_USER_WIDTH     => C_S_AXIS_USER_WIDTH,
      C_TRN_NP_FC             => C_TRN_NP_FC
      --C_M_AXI_AWUSER_WIDTH    => C_M_AXI_AWUSER_WIDTH,
      --C_M_AXI_WUSER_WIDTH     => C_M_AXI_WUSER_WIDTH
      --C_M_AXI_BUSER_WIDTH     => C_M_AXI_BUSER_WIDTH
      )
   port map(
      --AXI Global
      aclk                    => axi_aclk,
      reset                   => reset,
      --AXI Master Write Address Channel
      --m_axi_awid              => m_axi_awid,            --temporary
      m_axi_awaddr            => m_axi_awaddr,
      m_axi_awlen             => m_axi_awlen,
      m_axi_awsize            => m_axi_awsize,
      m_axi_awburst           => m_axi_awburst,
      m_axi_awprot            => m_axi_awprot,
      m_axi_awvalid           => m_axi_awvalid,
      m_axi_awready           => m_axi_awready,
      m_axi_awlock            => m_axi_awlock,
      m_axi_awcache           => m_axi_awcache,
      --m_axi_awuser     => m_axi_awuser,
      --AXI Master Write Data Channel
      m_axi_wdata             => m_axi_wdata,
      m_axi_wstrb             => m_axi_wstrb,
      m_axi_wlast             => m_axi_wlast,
      m_axi_wvalid            => m_axi_wvalid,
      m_axi_wready            => m_axi_wready,
      --m_axi_wuser      => m_axi_wuser,
      --AXI Master Write Response Channel
      m_axi_bresp             => m_axi_bresp,
      m_axi_bvalid            => m_axi_bvalid,
      m_axi_bready            => m_axi_bready,
      --m_axi_buser      => m_axi_buser,
      --Master Bridge Interrupt Strobes
      --master_int       => open,            --temporary
      MDE_int                 => MDE_int,
      MSE_int                 => MSE_int,
      MEP_int                 => MEP_int,
      --MLE_int                 => MLE_int,
      --MEC_int                 => MEC_int,
      --AXIS Write Completer Channel
      s_axis_cw_tdata         => s_axis_cw_tdata,
      s_axis_cw_tstrb         => s_axis_cw_tstrb,
      s_axis_cw_tlast         => s_axis_cw_tlast,
      s_axis_cw_tvalid        => s_axis_cw_tvalid,
      s_axis_cw_tready        => s_axis_cw_tready,
      s_axis_cw_tuser         => s_axis_cw_tuser,
      --AXI Master Read Address Channel
      --m_axi_arid              => m_axi_arid,
      m_axi_araddr            => m_axi_araddr,
      m_axi_arlen             => m_axi_arlen,
      m_axi_arsize            => m_axi_arsize,
      m_axi_arburst           => m_axi_arburst,
      m_axi_arprot            => m_axi_arprot,
      m_axi_arvalid           => m_axi_arvalid,
      m_axi_arready           => m_axi_arready,
      m_axi_arlock            => m_axi_arlock,
      m_axi_arcache           => m_axi_arcache,
    --m_axi_aruser     => m_axi_aruser,
    --AXI Master Read Data Channel
      m_axi_rdata             => m_axi_rdata,
      m_axi_rresp             => m_axi_rresp,
      m_axi_rlast             => m_axi_rlast,
      m_axi_rvalid            => m_axi_rvalid,
      m_axi_rready            => m_axi_rready,
    --m_axi_ruser      => m_axi_ruser,
    --AXIS Read Completer Channel
      s_axis_cr_tdata         => s_axis_cr_tdata,
      s_axis_cr_tstrb         => s_axis_cr_tstrb,
      s_axis_cr_tlast         => s_axis_cr_tlast,
      s_axis_cr_tvalid        => s_axis_cr_tvalid,
      s_axis_cr_tready        => s_axis_cr_tready,
      s_axis_cr_tuser         => s_axis_cr_tuser,
    --AXIS Completion Completer Channel
      m_axis_cc_tdata         => m_axis_cc_tdata,
      m_axis_cc_tstrb         => m_axis_cc_tstrb,
      m_axis_cc_tlast         => m_axis_cc_tlast,
      m_axis_cc_tvalid        => m_axis_cc_tvalid,
      m_axis_cc_tready        => m_axis_cc_tready,
      m_axis_cc_tuser         => m_axis_cc_tuser,
      --AXI Streaming Block Interface
      blk_lnk_up              => blk_lnk_up,
      blk_dcontrol            => blk_dcontrol,
      blk_bus_number          => blk_bus_number,
      blk_device_number       => blk_device_number,
      blk_function_number     => blk_function_number,
      --Internal Interface Ordering
      slwrreqpend             => slwrreqpendsig,
      slwrreqcomp             => slwrreqcompsig,
      wrreqpend               => wrreqpendsig,
      wrreqcomp               => wrreqcompsig,
      slv_write_idle          => sig_slv_write_idle,
      s_axi_awvalid           => sig_s_axi_awvalid,
      master_wr_idle          => sig_master_wr_idle,
      -- signals required for X7 NP credit return logic
      rdndreqpipeline         => rdndreqpipeline,
      rdreqpipeline           => rdreqpipeline,
      np_pkt_complete         => np_pkt_complete
      );

   comp_slave_bridge : entity axi_pcie_v2_9_14.slave_bridge
   generic map(
      --Family Generics
      C_FAMILY                      => C_FAMILY,
      C_S_AXI_ID_WIDTH              => C_S_AXI_ID_WIDTH,
      C_S_AXI_ADDR_WIDTH            => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH            => C_S_AXI_DATA_WIDTH,
      C_M_AXIS_DATA_WIDTH           => C_M_AXIS_DATA_WIDTH,
      C_COMP_TIMEOUT                => C_COMP_TIMEOUT,
      C_USER_CLK_FREQ               => C_USER_CLK_FREQ,
      C_USER_CLK2_DIV2              => C_USER_CLK2_DIV2,
      C_INCLUDE_RC                  => C_INCLUDE_RC,
      C_S_AXI_SUPPORTS_NARROW_BURST => C_S_AXI_SUPPORTS_NARROW_BURST,
      C_EP_LINK_PARTNER_RCB         => C_EP_LINK_PARTNER_RCB,
      C_AXIREAD_NUM                 => C_AXIREAD_NUM,   -- CR # 646225
      C_AXIBAR_NUM                  => C_AXIBAR_NUM,
      C_AXIBAR_0                    => C_AXIBAR_0,
      C_AXIBAR_AS_0                 => C_AXIBAR_AS_0,
      C_AXIBAR_AS_1                 => C_AXIBAR_AS_1,
      C_AXIBAR_AS_2                 => C_AXIBAR_AS_2,
      C_AXIBAR_AS_3                 => C_AXIBAR_AS_3,
      C_AXIBAR_AS_4                 => C_AXIBAR_AS_4,
      C_AXIBAR_AS_5                 => C_AXIBAR_AS_5,
      C_AXIBAR_HIGHADDR_0           => C_AXIBAR_HIGHADDR_0,
      C_AXIBAR_1                    => C_AXIBAR_1,
      C_AXIBAR_HIGHADDR_1           => C_AXIBAR_HIGHADDR_1,
      C_AXIBAR_2                    => C_AXIBAR_2,
      C_AXIBAR_HIGHADDR_2           => C_AXIBAR_HIGHADDR_2,
      C_AXIBAR_3                    => C_AXIBAR_3,
      C_AXIBAR_HIGHADDR_3           => C_AXIBAR_HIGHADDR_3,
      C_AXIBAR_4                    => C_AXIBAR_4,
      C_AXIBAR_HIGHADDR_4           => C_AXIBAR_HIGHADDR_4,
      C_AXIBAR_5                    => C_AXIBAR_5,
      C_AXIBAR_HIGHADDR_5           => C_AXIBAR_HIGHADDR_5,
      C_AXIBAR_CHK_SLV_ERR          => C_AXIBAR_CHK_SLV_ERR
   )
   port map(

      -- AXI Global
      s_axi_aclk              => axi_aclk,
      reset                   => reset,

      -- AXI Slave Write Address Channel
      s_axi_awid              => s_axi_awid,
      s_axi_awaddr            => s_axi_awaddr,
      s_axi_awregion          => s_axi_awregion,
      s_axi_awlen             => s_axi_awlen,
      s_axi_awsize            => s_axi_awsize,
      s_axi_awburst           => s_axi_awburst,
      s_axi_awvalid           => s_axi_awvalid,
      s_axi_awready           => s_axi_awready,

      -- AXI Slave Write Data Channel
      s_axi_wdata             => s_axi_wdata,
      s_axi_wstrb             => s_axi_wstrb,
      s_axi_wlast             => s_axi_wlast,
      s_axi_wvalid            => s_axi_wvalid,
      s_axi_wready            => s_axi_wready,

      -- AXI Slave Write Response Channel
      s_axi_bid               => s_axi_bid,
      s_axi_bresp             => s_axi_bresp,
      s_axi_bvalid            => s_axi_bvalid,
      s_axi_bready            => s_axi_bready,

      -- AXI Slave Read Address Channel
      s_axi_arid              => s_axi_arid,
      s_axi_araddr            => s_axi_araddr,
      s_axi_arregion          => s_axi_arregion,
      s_axi_arlen             => s_axi_arlen,
      s_axi_arsize            => s_axi_arsize,
      s_axi_arburst           => s_axi_arburst,
      s_axi_arvalid           => s_axi_arvalid,
      s_axi_arready           => s_axi_arready,

      -- AXI Slave Read Data Channel
      s_axi_rid               => s_axi_rid,
      s_axi_rdata             => s_axi_rdata,
      s_axi_rresp             => s_axi_rresp,
      s_axi_rlast             => s_axi_rlast,
      s_axi_rvalid            => s_axi_rvalid,
      s_axi_rready            => s_axi_rready,

      -- AXIS Write Requester Channel
      m_axis_rw_tdata         => m_axis_rw_tdata,
      m_axis_rw_tstrb         => m_axis_rw_tstrb,
      m_axis_rw_tlast         => m_axis_rw_tlast,
      m_axis_rw_tvalid        => m_axis_rw_tvalid,
      m_axis_rw_tready        => m_axis_rw_tready,

      -- AXIS Read Requester Channel
      m_axis_rr_tid           => m_axis_rr_tid,
      m_axis_rr_tdata         => m_axis_rr_tdata,
      m_axis_rr_tstrb         => m_axis_rr_tstrb,
      m_axis_rr_tlast         => m_axis_rr_tlast,
      m_axis_rr_tvalid        => m_axis_rr_tvalid,
      m_axis_rr_tready        => m_axis_rr_tready,

      -- AXIS Completion Requester Channel
      s_axis_rc_tdata         => s_axis_rc_tdata,
      s_axis_rc_tstrb         => s_axis_rc_tstrb,
      s_axis_rc_tlast         => s_axis_rc_tlast,
      s_axis_rc_tvalid        => s_axis_rc_tvalid,
      s_axis_rc_tready        => s_axis_rc_tready,

      -- AXI2PCIE translation vectors
      axibar2pciebar0         => axibar2pciebar0,
      axibar2pciebar1         => axibar2pciebar1,
      axibar2pciebar2         => axibar2pciebar2,
      axibar2pciebar3         => axibar2pciebar3,
      axibar2pciebar4         => axibar2pciebar4,
      axibar2pciebar5         => axibar2pciebar5,
      
      -- AXI-S Block Interface
      blk_lnk_up              => blk_lnk_up,
      blk_bus_number          => blk_bus_number,
      blk_device_number       => blk_device_number,
      blk_function_number     => blk_function_number,
      blk_command             => blk_command,
      blk_dcontrol            => blk_dcontrol,
      blk_lstatus             => blk_lstatus,
      np_cpl_pending          => np_cpl_pending,
      RP_bridge_en            => RP_bridge_en,

      -- Ordering signals
      --slrdready               => slrdready,
      --slcplready              => slcplready,
      --slrdsend                => slrdsend,
      --slcplsend               => slcplsend,
      pend_slv_wr_cnt         => slwrreqpendsig,
      cmpl_slv_wr_cnt         => slwrreqcompsig,
      wrreqpend               => wrreqpendsig,
      wrreqcomp               => wrreqcompsig,
      slv_write_idle          => sig_slv_write_idle,
      master_wr_idle          => sig_master_wr_idle,
      s_axi_awvalid_o         => sig_s_axi_awvalid,
      -- Slave Bridge Interrupt Strobes
      SUR                     => SUR_int,
      SUC                     => SUC_int,
      SCT                     => SCT_int,
      SEP                     => SEP_int,
      SCA                     => SCA_int,
      SIB                     => SIB_int,
      config_gen_req          => config_gen_req
   );

--clk_user_intr <= slave_int & master_int;

end architecture;


------------------------------------------------------------------------------------------------------------------------
--
--
--    File:       axi_pcie_msi_irq.vhd
--
--
--*--------------------------------------------------------------------------------------------------------------------*
--*                                                                                                                    *
--*      revision history:                                                                                             *
--*                                                                                                                    *
--*      31.10.2013  RE       - Initial revision                                                                       *
--*                                                                                                                    *
--*--------------------------------------------------------------------------------------------------------------------*


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_misc.ALL;
USE ieee.numeric_std.ALL;


PACKAGE axi_pcie_msi_irq_pkg IS

  COMPONENT axi_pcie_msi_irq
    GENERIC(
      g_data_width     : natural range 1 TO 64 := 32
			);
    PORT(
      COM_ICLK_I             : IN    std_logic;
      COM_CCLK_I             : IN    std_logic;
      COM_SYSRST_I           : IN    std_logic;
      
      MSI_MSG_RCVD_I         : IN    std_logic;
      MSI_IRQ_NUM_I          : IN    std_logic_vector(15 DOWNTO  0);
      
      MSI_IRQ_OVERFLOW_REG_O : OUT   std_logic_vector(g_data_width-1 DOWNTO  0);
      MSI_IRQ_UNDERRUN_REG_O : OUT   std_logic_vector(g_data_width-1 DOWNTO  0);
      
      IRQ_CLR_I              : IN    std_logic;
      IRQ_CLR_REG_I          : IN    std_logic_vector(g_data_width-1 DOWNTO  0);
      
      IRQ_STATUS_REG_O       : OUT   std_logic_vector(g_data_width-1 DOWNTO  0)
      );
  END COMPONENT axi_pcie_msi_irq;

END PACKAGE axi_pcie_msi_irq_pkg;


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;


ENTITY axi_pcie_msi_irq IS
  GENERIC(
    g_data_width : natural range 1 TO 64 := 32
    );
  PORT(
    COM_ICLK_I             : IN    std_logic;
    COM_CCLK_I             : IN    std_logic;
    COM_SYSRST_I           : IN    std_logic;
    
    MSI_MSG_RCVD_I         : IN    std_logic;
    MSI_IRQ_NUM_I          : IN    std_logic_vector(15 DOWNTO  0);
    
    MSI_IRQ_OVERFLOW_REG_O : OUT   std_logic_vector(g_data_width-1 DOWNTO  0);
    MSI_IRQ_UNDERRUN_REG_O : OUT   std_logic_vector(g_data_width-1 DOWNTO  0);
    
    IRQ_CLR_I              : IN    std_logic;
    IRQ_CLR_REG_I          : IN    std_logic_vector(g_data_width-1 DOWNTO  0);
    
    IRQ_STATUS_REG_O       : OUT   std_logic_vector(g_data_width-1 DOWNTO  0)
    );
END ENTITY axi_pcie_msi_irq;


ARCHITECTURE behavior OF axi_pcie_msi_irq IS

  CONSTANT c_data_width : natural range 1 TO 64 := g_data_width;
  
  SIGNAL s_msi_irq_line : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_msi_irq_num  : unsigned(15 DOWNTO  0);
  SIGNAL s_rst_cda      : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_rst_cda_1    : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_rst_cdb      : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_rst_cdb_1    : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_com_sysrst_1 : std_logic;
  SIGNAL s_com_sysrst   : std_logic;
  SIGNAL s_arst         : std_logic_vector(g_data_width-1 DOWNTO  0);
  
  SIGNAL s_msi_irq_pulse_cda : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_msi_irq_pulse_cdb : std_logic_vector(g_data_width-1 DOWNTO  0);
  
  TYPE t_std_logic_vector_2DW0 IS ARRAY (natural range <>) OF std_logic_vector( 2 DOWNTO  0);
  SIGNAL s_msi_irq_pulse_cda_dlyd : t_std_logic_vector_2DW0(g_data_width-1 DOWNTO  0);
  
  TYPE t_unsigned_vector_3DW0 IS ARRAY (natural range <>) OF unsigned( 3 DOWNTO  0);
  SIGNAL s_msi_irq_cnt : t_unsigned_vector_3DW0(g_data_width-1 DOWNTO  0);
  
  SIGNAL s_msi_irq_clr_pulse    : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_msi_irq_cnt_overflow : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_msi_irq_cnt_underrun : std_logic_vector(g_data_width-1 DOWNTO  0);
  SIGNAL s_msi_irq_status       : std_logic_vector(g_data_width-1 DOWNTO  0);
  
  
BEGIN

  s_msi_irq_num <= unsigned(MSI_IRQ_NUM_I);
  
  COM_SYSRST: PROCESS(COM_CCLK_I, COM_SYSRST_I)
  BEGIN
    IF (COM_SYSRST_I = '1') THEN
      s_com_sysrst_1 <= '1';
      s_com_sysrst   <= '1';
    ELSE
      IF rising_edge(COM_CCLK_I) THEN
        s_com_sysrst_1 <= '0';
        s_com_sysrst   <= s_com_sysrst_1;
      END IF;
    END IF;
  END PROCESS COM_SYSRST;
  
  
  G_MSI_IRQ_CLR: FOR i IN g_data_width-1 DOWNTO 0 GENERATE
    s_msi_irq_clr_pulse(i) <= IRQ_CLR_REG_I(i) AND IRQ_CLR_I;
  END GENERATE G_MSI_IRQ_CLR;
  
  
  G_MSI_IRQ_LINE: FOR i IN g_data_width-1 DOWNTO 0 GENERATE
  
    PROCESS(COM_ICLK_I)
    BEGIN
      IF rising_edge(COM_ICLK_I) THEN
        IF (MSI_MSG_RCVD_I = '1' AND
            s_msi_irq_num( 4 DOWNTO 0) = TO_UNSIGNED(i, 5)
           ) THEN
          s_msi_irq_line(i) <= '1';
        ELSE
          s_msi_irq_line(i) <= '0';
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE G_MSI_IRQ_LINE;
  
  
  G_MSI_IRQ_PACD: FOR i IN g_data_width-1 DOWNTO 0 GENERATE
    
    TFF: PROCESS(COM_ICLK_I, s_rst_cda(i))
    BEGIN
      IF rising_edge(COM_ICLK_I) THEN
        IF (s_rst_cda(i) = '1') THEN
          s_msi_irq_pulse_cda(i) <= '0';
        ELSE
          s_msi_irq_pulse_cda(i) <= s_msi_irq_pulse_cda(i) XOR s_msi_irq_line(i);
        END IF;
      END IF;
    END PROCESS TFF;
    
    DFF: PROCESS(COM_CCLK_I, s_rst_cdb(i))
    BEGIN
      IF rising_edge(COM_CCLK_I) THEN
        IF (s_rst_cdb(i) = '1') THEN
          s_msi_irq_pulse_cda_dlyd(i) <= (OTHERS => '0');
        ELSE
          s_msi_irq_pulse_cda_dlyd(i) <= s_msi_irq_pulse_cda_dlyd(i)(s_msi_irq_pulse_cda_dlyd(i)'high-1 DOWNTO  0) & s_msi_irq_pulse_cda(i);
        END IF;
      END IF;
    END PROCESS DFF;
    
    s_arst(i)              <= s_msi_irq_pulse_cda_dlyd(i)(s_msi_irq_pulse_cda_dlyd(i)'high) OR COM_SYSRST_I;
    s_msi_irq_pulse_cdb(i) <= s_msi_irq_pulse_cda_dlyd(i)(s_msi_irq_pulse_cda_dlyd(i)'high) XOR s_msi_irq_pulse_cda_dlyd(i)(s_msi_irq_pulse_cda_dlyd(i)'high-1);
    
    
    RST_TFF: PROCESS(COM_ICLK_I, s_arst(i))
    BEGIN
      IF (s_arst(i) = '1') THEN
        s_rst_cda_1(i) <= '1';
        s_rst_cda(i)   <= '1';
      ELSE
        IF rising_edge(COM_ICLK_I) THEN
          s_rst_cda_1(i) <= '0';
          s_rst_cda(i)   <= s_rst_cda_1(i);
        END IF;
      END IF;
    END PROCESS RST_TFF;
    
    RST_DFF: PROCESS(COM_CCLK_I, s_arst(i))
    BEGIN
      IF (s_arst(i) = '1') THEN
        s_rst_cdb_1(i) <= '1';
        s_rst_cdb(i)   <= '1';
      ELSE
        IF rising_edge(COM_CCLK_I) THEN
          s_rst_cdb_1(i) <= '0';
          s_rst_cdb(i)   <= s_rst_cdb_1(i);
        END IF;
      END IF;
    END PROCESS RST_DFF;
        
  END GENERATE G_MSI_IRQ_PACD;
  
  
  G_MSI_IRQ_CNT: FOR i IN g_data_width-1 DOWNTO  0 GENERATE
  
    MSI_IRQ_CNT: PROCESS(COM_CCLK_I, s_com_sysrst)
    BEGIN
      IF (s_com_sysrst = '1') THEN
        s_msi_irq_cnt(i)          <= to_unsigned(0, 4);
        s_msi_irq_cnt_overflow(i) <= '0';
        s_msi_irq_cnt_underrun(i) <= '0';
        s_msi_irq_status(i)       <= '0';
      ELSE
        IF rising_edge(COM_CCLK_I) THEN
          IF (s_msi_irq_pulse_cdb(i) = '1' AND s_msi_irq_clr_pulse(i) = '1') THEN
            s_msi_irq_cnt(i) <= s_msi_irq_cnt(i);
          ELSIF (s_msi_irq_pulse_cdb(i) = '1') THEN
            IF (s_msi_irq_cnt(i) < to_unsigned(15, 4)) THEN
              s_msi_irq_cnt(i)          <= s_msi_irq_cnt(i) + to_unsigned(1, 4);
              s_msi_irq_cnt_underrun(i) <= '0';
              s_msi_irq_status(i)       <= '1';
            ELSE
              s_msi_irq_cnt(i)          <= s_msi_irq_cnt(i);
              s_msi_irq_cnt_overflow(i) <= '1';
            END IF;
          ELSIF (s_msi_irq_clr_pulse(i) = '1') THEN
            IF (s_msi_irq_cnt(i) > to_unsigned(0, 4)) THEN
              s_msi_irq_cnt(i)          <= s_msi_irq_cnt(i) - to_unsigned(1, 4);
              s_msi_irq_cnt_overflow(i) <= '0';
              IF (s_msi_irq_cnt(i) = to_unsigned(1, 4)) THEN
                s_msi_irq_status(i) <= '0';
              ELSE
                s_msi_irq_status(i) <= s_msi_irq_status(i);
              END IF;
            ELSE
              s_msi_irq_cnt(i)          <= s_msi_irq_cnt(i);
              s_msi_irq_cnt_underrun(i) <= '1';
            END IF;
          END IF;
        END IF;
      END IF;
    END PROCESS MSI_IRQ_CNT;
    
    MSI_IRQ_OVERFLOW_REG_O(i) <= s_msi_irq_cnt_overflow(i);
    MSI_IRQ_UNDERRUN_REG_O(i) <= s_msi_irq_cnt_underrun(i);
    
  END GENERATE G_MSI_IRQ_CNT;
  
  
  IRQ_STATUS_REG_O <= s_msi_irq_status;
  
   
END ARCHITECTURE behavior;


-------------------------------------------------------------------------------
-- (c) Copyright 2020-2023 AMD, Inc. All rights reserved.
--
-- This file contains confidential and proprietary information
-- of AMD, Inc. and is protected under U.S. and 
-- international copyright and other intellectual property
-- laws.
--
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- AMD, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) AMD shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or AMD had been advised of the
-- possibility of the same.
--
-- CRITICAL APPLICATIONS
-- AMD products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of AMD products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
--
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
-- Filename:        axi_pcie.vhd
--
-- Description:     
--                  
-- This VHDL file is the HDL design file for the AXI PCIe bridge. 
--                   
-- Comments:
--                  
--                  
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--                axi_pcie.vhd
--
-------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.std_logic_misc.all;
--use ieee.std_logic_arith.conv_integer;
use ieee.std_logic_arith.conv_std_logic_vector;

library axi_pcie_v2_9_14;
use axi_pcie_v2_9_14.all;

--------------------------------------------------------------------------------
--Notes
--------------------------------------------------------------------------------



entity axi_pcie is
   generic(
      --Family Generics
      C_PCIE_BLK_LOCN               : string  := "0";
      C_XLNX_REF_BOARD              : string  := "NONE";
      C_FAMILY                      : string  := "virtex7";
      C_DEVICE                      : string  := "xc7k325t";
      C_SPEED                       : string  := "-1";
      C_INSTANCE                    : string  := "AXI_PCIe";
      C_S_AXI_ID_WIDTH              : integer := 4;
      -- C_M_AXI_THREAD_ID_WIDTH       : integer := 4;
      C_S_AXI_ADDR_WIDTH            : integer := 32;
      C_S_AXI_DATA_WIDTH            : integer := 32;
      C_M_AXI_ADDR_WIDTH            : integer := 32;
      C_M_AXI_DATA_WIDTH            : integer := 32;
    
      --PCIe Generics
      C_NO_OF_LANES                 : integer := 1;
      C_MAX_LINK_SPEED              : integer := 0;
                             -- 0 = 2.5 GT/s, 1 = 5.0 GT/s
      C_PCIE_USE_MODE               : string  := "1.0";
      C_DEVICE_ID                   : std_logic_vector := x"0000";
      C_VENDOR_ID                   : std_logic_vector := x"0000";
      C_CLASS_CODE                  : std_logic_vector := x"000000";
      C_REF_CLK_FREQ                : integer := 0;
                             --0 - 100 MHz, 1 - 125 MHz, 2 - 250 MHz
      PCIE_EXT_CLK                  : string:= "FALSE";
      EXT_PIPE_INTERFACE            : string:= "FALSE";
      PCIE_EXT_GT_COMMON            : string:= "FALSE";
      EXT_CH_GT_DRP                 : string:= "FALSE";
      SHARED_LOGIC_IN_CORE          : string:= "FALSE";
      TRANSCEIVER_CTRL_STATUS_PORTS : string:= "FALSE";
      AXI_ACLK_LOOPBACK             : string:= "FALSE";
      NO_SLV_ERR                    : string:= "FALSE";
      C_RP_BAR_HIDE                 : string:= "FALSE";
      C_TRN_NP_FC                   : string:= "FALSE";

      C_REV_ID                      : std_logic_vector := x"00";
      C_SUBSYSTEM_ID                : std_logic_vector := x"0000";
      C_SUBSYSTEM_VENDOR_ID         : std_logic_vector := x"0000";
      C_PCIE_CAP_SLOT_IMPLEMENTED   : integer := 0;
      C_SLOT_CLOCK_CONFIG           : string:= "TRUE";
      C_MSI_DECODE_ENABLE           : string:= "TRUE";
      C_NUM_MSI_REQ                 : integer := 0;
      C_INTERRUPT_PIN               : integer := 0;
      C_COMP_TIMEOUT                : integer := 0;
      C_INCLUDE_RC                  : integer := 0;
      C_S_AXI_SUPPORTS_NARROW_BURST : integer := 1;
      C_EP_LINK_PARTNER_RCB         : integer := 0;
      C_INCLUDE_BAROFFSET_REG       : integer := 1;
      C_BASEADDR                    : std_logic_vector := x"FFFF_FFFF";
      C_HIGHADDR                    : std_logic_vector := x"0000_0000";
      C_AXIBAR_NUM                  : integer := 6;
      C_AXIBAR2PCIEBAR_0            : std_logic_vector :=x"00000000";
      C_AXIBAR2PCIEBAR_1            : std_logic_vector :=x"00000000";
      C_AXIBAR2PCIEBAR_2            : std_logic_vector :=x"00000000";
      C_AXIBAR2PCIEBAR_3            : std_logic_vector :=x"00000000";
      C_AXIBAR2PCIEBAR_4            : std_logic_vector :=x"00000000";
      C_AXIBAR2PCIEBAR_5            : std_logic_vector :=x"00000000";
      C_AXIBAR_AS_0                 : integer := 0;
      C_AXIBAR_AS_1                 : integer := 0;
      C_AXIBAR_AS_2                 : integer := 0;
      C_AXIBAR_AS_3                 : integer := 0;
      C_AXIBAR_AS_4                 : integer := 0;
      C_AXIBAR_AS_5                 : integer := 0;
      C_AXIBAR_0                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_0           : std_logic_vector := x"0000_0000";
      C_AXIBAR_1                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_1           : std_logic_vector := x"0000_0000";
      C_AXIBAR_2                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_2           : std_logic_vector := x"0000_0000";
      C_AXIBAR_3                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_3           : std_logic_vector := x"0000_0000";
      C_AXIBAR_4                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_4           : std_logic_vector := x"0000_0000";
      C_AXIBAR_5                    : std_logic_vector := x"FFFF_FFFF";
      C_AXIBAR_HIGHADDR_5           : std_logic_vector := x"0000_0000";
      C_PCIEBAR_NUM                 : integer := 3;
      C_PCIEBAR_AS                  : integer := 1;
      C_PCIEBAR_LEN_0               : integer := 16;
      C_PCIEBAR2AXIBAR_0            : std_logic_vector(0 to 31) :=x"00000000";
      C_PCIEBAR2AXIBAR_0_SEC        : integer := 1;
      C_PCIEBAR_LEN_1               : integer := 16;
      C_PCIEBAR2AXIBAR_1            : std_logic_vector(0 to 31) :=x"00000000";
      C_PCIEBAR2AXIBAR_1_SEC        : integer := 1;
      C_PCIEBAR_LEN_2               : integer := 16;
      C_PCIEBAR2AXIBAR_2            : std_logic_vector(0 to 31) :=x"00000000";
      C_PCIEBAR2AXIBAR_2_SEC        : integer := 1;
      ENABLE_JTAG_DBG               : string := "FALSE";
      REDUCE_OOB_FREQ               : string := "FALSE";
      C_INT_FIFO_DEPTH              : integer := 0;
      C_AXIBAR_CHK_SLV_ERR          : string := "FALSE"
   );
   port(
      -- AXI Global
      axi_aclk                : in  std_logic; -- AXI clock
      axi_aresetn             : in  std_logic; -- AXI active low synchronous reset
      axi_aclk_out            : out std_logic; -- PCIe clock for AXI clock
      axi_ctl_aclk            : in  std_logic; -- AXI LITE clock
      axi_ctl_aclk_out        : out std_logic; -- PCIe clock for AXI LITE clock
      mmcm_lock               : out std_logic := '1'; -- MMCM lock signal output
      user_link_up            : out std_logic; -- user linkup signal output
      interrupt_out           : out std_logic; -- active high interrupt out
      INTX_MSI_Request        : in  std_logic; -- Legacy interrupt/initiate MSI (Endpoint only)
      INTX_MSI_Grant          : out std_logic; -- Legacy interrupt/MSI Grant signal (Endpoint only)
      MSI_enable              : out std_logic; -- 1 = MSI, 0 = INTX
      MSI_Vector_Num          : in  std_logic_vector(4 downto 0);
      MSI_Vector_Width        : out std_logic_vector(2 downto 0);

      -- AXI Slave Write Address Channel
      s_axi_awid              : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_awaddr            : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_awregion          : in  std_logic_vector(3 downto 0);
      s_axi_awlen             : in  std_logic_vector(7 downto 0);
      s_axi_awsize            : in  std_logic_vector(2 downto 0);
      s_axi_awburst           : in  std_logic_vector(1 downto 0);
      s_axi_awvalid           : in  std_logic;
      s_axi_awready           : out std_logic;

      -- AXI Slave Write Data Channel
      s_axi_wdata             : in  std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_wstrb             : in  std_logic_vector(C_S_AXI_DATA_WIDTH/8-1 downto 0);
      s_axi_wlast             : in  std_logic;
      s_axi_wvalid            : in  std_logic;
      s_axi_wready            : out std_logic;

      -- AXI Slave Write Response Channel
      s_axi_bid               : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_bresp             : out std_logic_vector(1 downto 0);
      s_axi_bvalid            : out std_logic;
      s_axi_bready            : in  std_logic;

      -- AXI Slave Read Address Channel
      s_axi_arid              : in  std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_araddr            : in  std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
      s_axi_arregion          : in  std_logic_vector(3 downto 0);
      s_axi_arlen             : in  std_logic_vector(7 downto 0);
      s_axi_arsize            : in  std_logic_vector(2 downto 0);
      s_axi_arburst           : in  std_logic_vector(1 downto 0);
      s_axi_arvalid           : in  std_logic;
      s_axi_arready           : out std_logic;

      -- AXI Slave Read Data Channel
      s_axi_rid               : out std_logic_vector(C_S_AXI_ID_WIDTH-1 downto 0);
      s_axi_rdata             : out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
      s_axi_rresp             : out std_logic_vector(1 downto 0);
      s_axi_rlast             : out std_logic;
      s_axi_rvalid            : out std_logic;
      s_axi_rready            : in  std_logic;

      -- AXI Master Write Address Channel
      m_axi_awaddr            : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
      m_axi_awlen             : out std_logic_vector(7 downto 0);
      m_axi_awsize            : out std_logic_vector(2 downto 0);
      m_axi_awburst           : out std_logic_vector(1 downto 0);
      m_axi_awprot            : out std_logic_vector(2 downto 0);
      m_axi_awvalid           : out std_logic;
      m_axi_awready           : in  std_logic;
      --m_axi_awid              : out std_logic_vector(C_M_AXI_THREAD_ID_WIDTH-1 downto 0);
      m_axi_awlock            : out std_logic;
      m_axi_awcache           : out std_logic_vector(3 downto 0);

      -- AXI Master Write Data Channel
      m_axi_wdata             : out std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
      m_axi_wstrb             : out std_logic_vector(C_M_AXI_DATA_WIDTH/8-1 downto 0);
      m_axi_wlast             : out std_logic;
      m_axi_wvalid            : out std_logic;
      m_axi_wready            : in  std_logic;

      -- AXI Master Write Response Channel
      m_axi_bresp             : in  std_logic_vector(1 downto 0);
      m_axi_bvalid            : in  std_logic;
      m_axi_bready            : out std_logic;

      -- AXI Master Read Address Channel
      --m_axi_arid              : out std_logic_vector(C_M_AXI_THREAD_ID_WIDTH-1 downto 0);
      m_axi_araddr            : out std_logic_vector(C_M_AXI_ADDR_WIDTH-1 downto 0);
      m_axi_arlen             : out std_logic_vector(7 downto 0);
      m_axi_arsize            : out std_logic_vector(2 downto 0);
      m_axi_arburst           : out std_logic_vector(1 downto 0);
      m_axi_arprot            : out std_logic_vector(2 downto 0);
      m_axi_arvalid           : out std_logic;
      m_axi_arready           : in  std_logic;
      m_axi_arlock            : out std_logic;
      m_axi_arcache           : out std_logic_vector(3 downto 0);

      -- AXI Master Read Data Channel
      m_axi_rdata             : in  std_logic_vector(C_M_AXI_DATA_WIDTH-1 downto 0);
      m_axi_rresp             : in  std_logic_vector(1 downto 0);
      m_axi_rlast             : in  std_logic;
      m_axi_rvalid            : in  std_logic;
      m_axi_rready            : out std_logic;

      -- PCI Express (pci_exp) Interface
      -- Tx
      pci_exp_txp             : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
      pci_exp_txn             : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
      -- Rx
      pci_exp_rxp             : in  std_logic_vector(C_NO_OF_LANES-1 downto 0);
      pci_exp_rxn             : in  std_logic_vector(C_NO_OF_LANES-1 downto 0);
      REFCLK                  : in  std_logic;
      

      -- AXI -Lite Interface - CFG Block
      s_axi_ctl_awaddr        : in  std_logic_vector(31 downto 0); -- AXI Lite Write address
      s_axi_ctl_awvalid       : in  std_logic;                     -- AXI Lite Write Address Valid
      s_axi_ctl_awready       : out std_logic;                     -- AXI Lite Write Address Core ready
      s_axi_ctl_wdata         : in  std_logic_vector(31 downto 0); -- AXI Lite Write Data
      s_axi_ctl_wstrb         : in  std_logic_vector(3 downto 0);  -- AXI Lite Write Data strobe
      s_axi_ctl_wvalid        : in  std_logic;                     -- AXI Lite Write data Valid
      s_axi_ctl_wready        : out std_logic;                     -- AXI Lite Write Data Core ready
      s_axi_ctl_bresp         : out std_logic_vector(1 downto 0);  -- AXI Lite Write Data strobe
      s_axi_ctl_bvalid        : out std_logic;                     -- AXI Lite Write data Valid
      s_axi_ctl_bready        : in  std_logic;                     -- AXI Lite Write Data Core ready

      s_axi_ctl_araddr        : in  std_logic_vector(31 downto 0); -- AXI Lite Read address
      s_axi_ctl_arvalid       : in  std_logic;                     -- AXI Lite Read Address Valid
      s_axi_ctl_arready       : out std_logic;                     -- AXI Lite Read Address Core ready
      s_axi_ctl_rdata         : out std_logic_vector(31 downto 0); -- AXI Lite Read Data
      s_axi_ctl_rresp         : out std_logic_vector(1 downto 0);  -- AXI Lite Read Data strobe
      s_axi_ctl_rvalid        : out std_logic;                     -- AXI Lite Read data Valid
      s_axi_ctl_rready        : in  std_logic;                     -- AXI Lite Read Data Core ready
qpll_drp_crscode      : in std_logic_vector(11 downto 0);
 qpll_drp_fsm          : in std_logic_vector(17 downto 0);
 qpll_drp_done         : in std_logic_vector(1 downto 0);
 qpll_drp_reset        : in std_logic_vector(1 downto 0);
 qpll_qplllock         : in std_logic_vector(1 downto 0);
 qpll_qplloutclk       : in std_logic_vector(1 downto 0);
 qpll_qplloutrefclk    : in std_logic_vector(1 downto 0);
  qpll_qplld    : out std_logic_vector(1 downto 0)        ;
  qpll_qpllreset: out std_logic_vector(1 downto 0)    ;
  qpll_drp_clk: out std_logic_vector(1 downto 0)    ;
  qpll_drp_rst_n: out std_logic_vector(1 downto 0)    ;
  qpll_drp_ovrd: out std_logic_vector(1 downto 0)    ;
  qpll_drp_gen3: out std_logic_vector(1 downto 0)    ;
  qpll_drp_start: out std_logic_vector(1 downto 0)    ;

  pipe_txprbssel               :in std_logic_vector(2 downto 0);
  pipe_rxprbssel               :in std_logic_vector(2 downto 0);
  pipe_txprbsforceerr  :in std_logic;
  pipe_rxprbscntreset  :in std_logic;
  pipe_loopback                :in std_logic_vector(2 downto 0);
  pipe_txinhibit               :in std_logic_vector(C_NO_OF_LANES-1 downto 0);

  pipe_rxprbserr : out std_logic_vector(C_NO_OF_LANES-1 downto 0);


  pipe_rst_fsm         :out std_logic_vector(4 downto 0);
  pipe_qrst_fsm        :out std_logic_vector(11 downto 0);
  pipe_rate_fsm        :out std_logic_vector((C_NO_OF_LANES*5)-1 downto 0);
  pipe_sync_fsm_tx     :out std_logic_vector((C_NO_OF_LANES*6)-1 downto 0);
  pipe_sync_fsm_rx     :out std_logic_vector((C_NO_OF_LANES*7)-1 downto 0);
  pipe_drp_fsm         :out std_logic_vector((C_NO_OF_LANES*7)-1 downto 0);

  pipe_rst_idle        :out std_logic;
  pipe_qrst_idle       :out std_logic;
  pipe_rate_idle       :out std_logic;
  pipe_eyescandataerror	:out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_rxstatus : out std_logic_vector((C_NO_OF_LANES*3)-1 downto 0);    
  pipe_dmonitorout : out std_logic_vector((C_NO_OF_LANES*15)-1 downto 0);

 pipe_cpll_lock          : out std_logic_vector(C_NO_OF_LANES-1 downto 0); 
 pipe_qpll_lock          : out std_logic_vector(((C_NO_OF_LANES/8)+1)-1 downto 0); 
 pipe_rxpmaresetdone     : out std_logic_vector(C_NO_OF_LANES-1 downto 0);  
 pipe_rxbufstatus        : out std_logic_vector((C_NO_OF_LANES*3)-1 downto 0);     
 pipe_txphaligndone      : out std_logic_vector(C_NO_OF_LANES-1 downto 0);   
 pipe_txphinitdone       : out std_logic_vector(C_NO_OF_LANES-1 downto 0);      
 pipe_txdlysresetdone    : out std_logic_vector(C_NO_OF_LANES-1 downto 0);    
 pipe_rxphaligndone      : out std_logic_vector(C_NO_OF_LANES-1 downto 0);     
 pipe_rxdlysresetdone    : out std_logic_vector(C_NO_OF_LANES-1 downto 0);      
 pipe_rxsyncdone         : out std_logic_vector(C_NO_OF_LANES-1 downto 0);      
 pipe_rxdisperr          : out std_logic_vector((C_NO_OF_LANES*8)-1 downto 0);     
 pipe_rxnotintable       : out std_logic_vector((C_NO_OF_LANES*8)-1 downto 0);     
 pipe_rxcommadet         : out std_logic_vector(C_NO_OF_LANES-1 downto 0);   

  gt_ch_drp_rdy        :out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_0 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_1 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_2 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_3 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_4 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_5 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_6 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_7 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_8 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug_9 : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
  pipe_debug   :out std_logic_vector(31 downto 0);

 common_commands_in:in std_logic_vector(11 downto 0); 	
 pipe_rx_0_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_1_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_2_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_3_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_4_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_5_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_6_sigs	   :in std_logic_vector(24 downto 0);     
 pipe_rx_7_sigs	   :in std_logic_vector(24 downto 0);     
                          
 common_commands_out:out std_logic_vector(11 downto 0);	
 pipe_tx_0_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_1_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_2_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_3_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_4_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_5_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_6_sigs	    :out std_logic_vector(24 downto 0);    
 pipe_tx_7_sigs	    :out std_logic_vector(24 downto 0);    

 int_pclk_out_slave	: out std_logic;	 
 int_rxusrclk_out    	: out std_logic;   	
 int_dclk_out        	: out std_logic;   	
 int_userclk1_out    	: out std_logic;   	
 int_userclk2_out    	: out std_logic;   	
 int_oobclk_out      	: out std_logic;   	
 int_mmcm_lock_out   	: out std_logic;   	
 int_qplllock_out	: out std_logic_vector(1 downto 0);	
 int_qplloutclk_out	: out std_logic_vector(1 downto 0);	
 int_qplloutrefclk_out	: out std_logic_vector(1 downto 0);	
 int_rxoutclk_out 	: out std_logic_vector(C_NO_OF_LANES-1 downto 0);	      
 int_pclk_sel_slave	: in std_logic_vector(C_NO_OF_LANES-1 downto 0);	

     -------------Channel DRP---------------------------------
  ext_ch_gt_drpclk      : out std_logic;
  ext_ch_gt_drpaddr     : in std_logic_vector((C_NO_OF_LANES*9)-1 downto 0);
  ext_ch_gt_drpen       : in std_logic_vector(C_NO_OF_LANES-1 downto 0);
  ext_ch_gt_drpdi       : in std_logic_vector((C_NO_OF_LANES*16)-1 downto 0);
  ext_ch_gt_drpwe       : in std_logic_vector(C_NO_OF_LANES-1 downto 0);

  ext_ch_gt_drpdo      : out std_logic_vector((C_NO_OF_LANES*16)-1 downto 0);
  ext_ch_gt_drprdy     : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
      clk_fab_refclk                           : in std_logic_vector(C_NO_OF_LANES-1 downto 0);
      clk_pclk                                 : in std_logic;
      clk_rxusrclk                             : in std_logic;
      clk_dclk                                 : in std_logic;
      clk_userclk1                             : in std_logic;
      clk_userclk2                             : in std_logic;
      clk_oobclk_in                            : in std_logic;
      clk_mmcm_lock                            : in std_logic;
      clk_txoutclk                             : out std_logic;
      clk_rxoutclk                             : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
      clk_pclk_sel                             : out std_logic_vector(C_NO_OF_LANES-1 downto 0);
      pipe_mmcm_rst_n                          : in std_logic;
      clk_gen3                                 : out std_logic
   );

end axi_pcie;

architecture structure of axi_pcie is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of structure : architecture is "yes";


-------------------------------------------------------------------------------

  -- Copied function "to_string" from MicroBlaze v8.30a
  
  -----------------------------------------------------------------------------
  -- Converts an integer to a decimal string
  -----------------------------------------------------------------------------
  function To_String(from : integer) return string is
  begin
    return integer'image(from);
  end function To_String;

  -----------------------------------------------------------------------------
  -- Converts a std_logic_vector to a hexadecimal string with leading "0x"
  -----------------------------------------------------------------------------
  function To_String(from : std_logic_vector) return String is
    type INT_TO_CHAR_TYPE is array (integer range 0 to 15) of character;
    constant INT_TO_STRHEX_TABLE : INT_TO_CHAR_TYPE :=
      ('0','1','2','3','4','5','6','7','8','9','A','B','C','D','E','F');

    variable value   : unsigned(0 to ((from'length + 3) / 4) * 4 - 1) := (others => '0');
    variable result  : string(1 to value'length / 4);
    variable v_index : integer := value'high;
    variable r_index : integer := result'high;
  begin
    value(value'high - from'length + 1 to value'high) := unsigned(from);
    while r_index > 0 loop
      result(r_index) := INT_TO_STRHEX_TABLE(to_integer(value(v_index - 3 to v_index)));
      v_index := v_index - 4;
      r_index := r_index - 1;
    end loop;
    return "0x" & result;
  end function To_String;


-------------------------------------------------------------------------------



  constant C_CORE_GENERATION_INFO : string := C_INSTANCE & ",AXI_PCIe,{"
      & "c_instance="                      & C_INSTANCE
      & ",c_family="                       & C_FAMILY
      & ",c_s_axi_id_width="               & to_string(C_S_AXI_ID_WIDTH)
      & ",c_s_axi_data_width="             & to_string(C_S_AXI_DATA_WIDTH)
      & ",c_m_axi_data_width="             & to_string(C_M_AXI_DATA_WIDTH)
      & ",c_no_of_lanes="                  & to_string(C_NO_OF_LANES)
      & ",c_max_link_speed="               & to_string(C_MAX_LINK_SPEED)
      & ",c_ref_clk_freq="                 & to_string(C_REF_CLK_FREQ)
      & ",c_pcie_cap_slot_implemented="   & to_string(C_PCIE_CAP_SLOT_IMPLEMENTED)
      & ",c_num_msi_req ="                 & to_string(C_NUM_MSI_REQ)
      & ",c_interrupt_pin="                & to_string(C_INTERRUPT_PIN)
      & ",c_include_rc="                   & to_string(C_INCLUDE_RC)
      & ",c_s_axi_supports_narrow_burst="  & to_string(C_S_AXI_SUPPORTS_NARROW_BURST)
      & ",c_include_baroffset_reg="      & to_string(C_INCLUDE_BAROFFSET_REG)
      & ",c_axibar_num="                   & to_string(C_AXIBAR_NUM)
      & ",c_pciebar_num="                 & to_string(C_PCIEBAR_NUM)
      & "}";

  attribute CORE_GENERATION_INFO : string;
  attribute CORE_GENERATION_INFO of structure : architecture is C_CORE_GENERATION_INFO;

-------------------------------------------------------------------------------

   function Conv_to_String(BINARY_INTEGER : integer) return string is
      begin
         if(BINARY_INTEGER = 0) then
            return("FALSE");
         else
            return("TRUE");
         end if;
   end function;
   function Conv_to_String_Inv(BINARY_INTEGER : integer) return string is
      begin
         if(BINARY_INTEGER = 1) then
            return("FALSE");
         else
            return("TRUE");
         end if;
   end function;
   function String_Inv(STRING_VAL : string) return string is
      begin
         if(STRING_VAL = "TRUE") then
            return("FALSE");
         else
            return("TRUE");
         end if;
   end function;

  constant CON_PCIE_CAP_SLOT_IMPLEMENTED : string := Conv_to_String(C_PCIE_CAP_SLOT_IMPLEMENTED);
  constant ROOT_PORT : string := Conv_to_String(C_INCLUDE_RC);
  constant UPSTREAM_FACING : string := Conv_to_String(1-C_INCLUDE_RC);
  constant VSEC_CAP_LAST : string := Conv_to_String(1-C_INCLUDE_BAROFFSET_REG);
  constant PCIE_ASYNC_EN : string := String_Inv(C_SLOT_CLOCK_CONFIG);
  
  
  
-------------------------------------------------------------------------------
-- prefetch_config
-- This function configures PCIBAR_PREFETCH parmameters
-------------------------------------------------------------------------------

--function prefetch_config(pcibar_as, use_prefetch_from_pkg, pcibar_prefetch : integer) return integer is
--   variable var_out : integer;
--   begin
--      if(use_prefetch_from_pkg=0) then
--         var_out := pcibar_as;
--      else
--         var_out := pcibar_prefetch;
--      end if;
--   return(var_out);
--end function;

-------------------------------------------------------------------------------
-- Function func_invert
-- This function takes in a SLV, inverts all bits in the vector and returns
-- a SLV
-------------------------------------------------------------------------------
  function func_invert(in_vec : std_logic_vector(63 downto 0)) return std_logic_vector is
    variable var_out : std_logic_vector(63 downto 0);
      begin
        for i in 0 to 63 loop
          var_out(i):=not in_vec(i);
        end loop;
      return(var_out);
  end function;

-------------------------------------------------------------------------------
-- pcibar_config
-- This function configures the PCIBARs
-------------------------------------------------------------------------------

  constant PCIBAR_PREFETCH_0  : integer := C_PCIEBAR_AS;  --prefetch_config(C_PCIEBAR_AS, 0, 0);
  constant PCIBAR_PREFETCH_1  : integer := C_PCIEBAR_AS;  --prefetch_config(C_PCIEBAR_AS, 0, 0);
  constant PCIBAR_PREFETCH_2  : integer := C_PCIEBAR_AS;  --prefetch_config(C_PCIEBAR_AS, 0, 0);

  function pcibar_config(pcibar_prefetch_32, pcibar_prefetch_64, pcibar_as, pcibar_len_32, pcibar_len_64, pcibar_en, pcibar_num_32, pcibar_num_64 : integer) return std_logic_vector is
     variable var_out : std_logic_vector(63 downto 0);
     begin
        if(pcibar_as=1) then -- 64 bit BARs
           if(pcibar_num_64<pcibar_en) then
              if(pcibar_prefetch_64=1) then
                 if (pcibar_len_64 = 32) then
                   var_out := x"FFFF_FFFF_0000_0000" + x"C";
                 elsif (pcibar_len_64 = 31) then
                   var_out := x"FFFF_FFFF_8000_0000" + x"C";
                 else
                   var_out := func_invert(conv_std_logic_vector(((2**pcibar_len_64)-1),64))+x"C";
                 end if;
              else
                 assert FALSE
                 report "INVALID BAR: 64 bit, non-prefetch NOT ALLOWED"
                 severity Warning;
              end if;
           else
              var_out:= (others=>'0');
           end if;
        else               -- 32 bit BARs
           if(pcibar_num_32<pcibar_en) then
              if(pcibar_prefetch_32=1) then
                 assert FALSE
                 report "INVALID BAR: 32 bit, prefetch NOT ALLOWED"
                 severity Warning;
              else
                 if(pcibar_num_32=1) then
                   if (pcibar_len_32 = 32) then
                     var_out := x"0000_0000"+x"0"&x"0000_0000";
                   elsif (pcibar_len_32 = 31) then
                     var_out := x"8000_0000"+x"0"&x"0000_0000";
                   else
                     var_out := func_invert(conv_std_logic_vector(((2**pcibar_len_32)-1),64))(31 downto 0)+x"0"&x"0000_0000";
                   end if;
                 else
                   if (pcibar_len_32 = 32) then
                     var_out := x"0000_0000"&x"0000_0000"+x"0";
                   elsif (pcibar_len_32 = 31) then
                     var_out := x"0000_0000"&x"8000_0000"+x"0";
                   else
                     var_out := x"0000_0000"&func_invert(conv_std_logic_vector(((2**pcibar_len_32)-1),64))(31 downto 0)+x"0";
                   end if;
                 end if;
              end if;
           else
              var_out := (others=>'0');
           end if;
        end if;
     return(var_out);
  end function;

  --------------------------------------------------------------------------------

  function group_7series_family (C_FAMILY : string) return string is
    begin
      if (C_FAMILY = "kintex7" or C_FAMILY = "virtex7" or C_FAMILY = "artix7" or C_FAMILY = "zynq") then
        return ("7series");
      else
        return (C_FAMILY);
      end if;
  end function;

  --------------------------------------------------------------------------------
  -- purpose: Assign the value to depending on the device port type 
  function get_dll_link_active_report_cap (
    constant dev_port : integer)
      return string is
   begin  -- get_dll_link_active_report_cap 
     if (dev_port = 1) then 
        return ("TRUE");
     else 
        return ("FALSE");
     end if; 
   end get_dll_link_active_report_cap;

  -- Added to find derivative of all FPGA architectures.
  -- For example, "virtex6l" will return "virtex6" (so correct V6 PCIe block is instantiated)
--  constant C_FAMILY_DER           : string := get_root_family (C_FAMILY);

  -- Added to group together 7-series FPGA architectures.
  constant C_FAMILY_I         : string := "7series";
  --constant C_FAMILY_I         : string := group_7series_family (C_FAMILY_DER);

  constant C_S_AXIS_DATA_WIDTH          : integer := C_S_AXI_DATA_WIDTH;
  constant C_M_AXIS_DATA_WIDTH          : integer := C_M_AXI_DATA_WIDTH;
  constant C_S_AXIS_USER_WIDTH          : integer := 22;
  constant NUM_OF_INTERRUPTS            : integer := 9;
  constant ZEROS                        : std_logic_vector(7 downto 0):= "00000000";
  constant BASEADDR_i                   : std_logic_vector(31 downto 0):= C_BASEADDR;
  constant BASEADDR_U                   : std_logic_vector(15 downto 0):= BASEADDR_i(31 downto 16);
  constant BASEADDR_L                   : std_logic_vector(15 downto 0):= BASEADDR_i(15 downto 0);
  constant HIGHADDR_i                   : std_logic_vector(31 downto 0):= C_HIGHADDR;
  constant HIGHADDR_U                   : std_logic_vector(15 downto 0):= HIGHADDR_i(31 downto 16);
  constant HIGHADDR_L                   : std_logic_vector(15 downto 0):= HIGHADDR_i(15 downto 0);
  constant PCIE_GENERIC                 : integer := conv_integer("010001101111") + (128*C_INTERRUPT_PIN);
  constant C_PL_FAST_TRAIN              : string := "FALSE"; --default hardware is not fast train
  constant LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP_LOCAL : string := get_dll_link_active_report_cap (C_INCLUDE_RC);
  constant MODELSIM                     : boolean := false --sim is always fast train
-- synthesis translate_off
       or true
-- synthesis translate_on
  ;

  function Fast_Train_Conv(MODELSIM : boolean; C_PL_FAST_TRAIN : string) return string is
    begin
      if(MODELSIM) then
        return("TRUE");
      else
-- coverage off
        return(C_PL_FAST_TRAIN);
-- coverage on
      end if;
  end function;

  constant C_PL_FAST_TRAIN_LOCAL : string := Fast_Train_Conv(MODELSIM, C_PL_FAST_TRAIN);
  constant BAR0_i  : std_logic_vector(31 downto 0):= pcibar_config(PCIBAR_PREFETCH_0, PCIBAR_PREFETCH_0, C_PCIEBAR_AS, C_PCIEBAR_LEN_0, C_PCIEBAR_LEN_0, C_PCIEBAR_NUM, 0, 0)(31 downto 0);
  constant BAR0_U  : std_logic_vector(15 downto 0):=BAR0_i(31 downto 16);
  constant BAR0_L  : std_logic_vector(15 downto 0):=BAR0_i(15 downto 0);
  constant BAR1_i  : std_logic_vector(31 downto 0):= pcibar_config(PCIBAR_PREFETCH_1, PCIBAR_PREFETCH_0, C_PCIEBAR_AS, C_PCIEBAR_LEN_1, C_PCIEBAR_LEN_0, C_PCIEBAR_NUM, 1, 0)(63 downto 32);
  constant BAR1_U  : std_logic_vector(15 downto 0):=BAR1_i(31 downto 16);
  constant BAR1_L  : std_logic_vector(15 downto 0):=BAR1_i(15 downto 0);
  constant BAR2_i  : std_logic_vector(31 downto 0):= pcibar_config(PCIBAR_PREFETCH_2, PCIBAR_PREFETCH_1, C_PCIEBAR_AS, C_PCIEBAR_LEN_2, C_PCIEBAR_LEN_1, C_PCIEBAR_NUM, 2, 1)(31 downto 0);
  constant BAR2_U_EP  : std_logic_vector(15 downto 0):=BAR2_i(31 downto 16);
  constant BAR2_L_EP  : std_logic_vector(15 downto 0):=BAR2_i(15 downto 0);
  constant BAR3_i  : std_logic_vector(31 downto 0):= pcibar_config(PCIBAR_PREFETCH_2, PCIBAR_PREFETCH_1, C_PCIEBAR_AS, C_PCIEBAR_LEN_2, C_PCIEBAR_LEN_1, C_PCIEBAR_NUM, 3, 1)(63 downto 32);
  constant BAR3_U_EP  : std_logic_vector(15 downto 0):=BAR3_i(31 downto 16);
  constant BAR3_L_EP  : std_logic_vector(15 downto 0):=BAR3_i(15 downto 0);
  constant BAR4_i  : std_logic_vector(31 downto 0):= pcibar_config(PCIBAR_PREFETCH_2, PCIBAR_PREFETCH_2, C_PCIEBAR_AS, C_PCIEBAR_LEN_2, C_PCIEBAR_LEN_2, C_PCIEBAR_NUM, 4, 2)(31 downto 0);
  constant BAR4_U_EP  : std_logic_vector(15 downto 0):=BAR4_i(31 downto 16);
  constant BAR4_L_EP  : std_logic_vector(15 downto 0):=BAR4_i(15 downto 0);
  constant BAR5_i  : std_logic_vector(31 downto 0):= pcibar_config(PCIBAR_PREFETCH_2, PCIBAR_PREFETCH_2, C_PCIEBAR_AS, C_PCIEBAR_LEN_2, C_PCIEBAR_LEN_2, C_PCIEBAR_NUM, 5, 2)(63 downto 32);
  constant BAR5_U_EP  : std_logic_vector(15 downto 0):=BAR5_i(31 downto 16);
  constant BAR5_L_EP  : std_logic_vector(15 downto 0):=BAR5_i(15 downto 0);
  --Fixed for V6 RP configuration
  constant BAR2_U_RP      : std_logic_vector(15 downto 0):=x"00ff";
  constant BAR2_L_RP      : std_logic_vector(15 downto 0):=x"ffff";
  constant BAR3_U_RP      : std_logic_vector(15 downto 0):=x"ffff";
  constant BAR3_L_RP      : std_logic_vector(15 downto 0):=x"f1f1";
  constant BAR4_U_RP      : std_logic_vector(15 downto 0):=x"fff0";
  constant BAR4_L_RP      : std_logic_vector(15 downto 0):=x"fff0";
  constant BAR5_U_RP      : std_logic_vector(15 downto 0):=x"0000";
  constant BAR5_L_RP      : std_logic_vector(15 downto 0):=x"0000";

-- coverage off

  --------------------------------------------------------------------------------

  function rp_bars_mux(C_INCLUDE_RC : integer; EP_BAR, RP_BAR : std_logic_vector) return std_logic_vector is
    begin
      if(C_INCLUDE_RC = 0) then
        return(EP_BAR);
      else
        return(RP_BAR);
      end if;
  end function;

  constant BAR2_U             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR2_U_EP, BAR2_U_RP);
  constant BAR2_L             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR2_L_EP, BAR2_L_RP);
  constant BAR3_U             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR3_U_EP, BAR3_U_RP);
  constant BAR3_L             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR3_L_EP, BAR3_L_RP);
  constant BAR4_U             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR4_U_EP, BAR4_U_RP);
  constant BAR4_L             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR4_L_EP, BAR4_L_RP);
  constant BAR5_U             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR5_U_EP, BAR5_U_RP);
  constant BAR5_L             : std_logic_vector  := rp_bars_mux(C_INCLUDE_RC, BAR5_L_EP, BAR5_L_RP);



  --------------------------------------------------------------------------------

  function set_pcie_use_mode (C_PCIE_USE_MODE : string) return string is
    begin
      -- Make sure C_PCI_USE_MODE = 3.0 for GES K7 GT wrappers in Zynq.  
      --if (C_FAMILY = "zynq") then
      --  return ("3.0");
      --else
        return (C_PCIE_USE_MODE);
      --end if;
  end function;

  constant PCIE_USE_MODE : string := set_pcie_use_mode (C_PCIE_USE_MODE);

  --------------------------------------------------------------------------------

  --------------------------------------------------------------------------------

  function set_pcie_gt_device (C_FAMILY : string) return string is
    begin
      -- Make sure  PCIE_GT_DEVICE = GTP for A7 GT wrappers.  
      if (C_FAMILY = "artix7" or (C_FAMILY = "zynq" and (C_DEVICE = "xc7z015" or C_DEVICE = "xc7z015i" or C_DEVICE = "xc7z012s"))) then
        return ("GTP");
      else
        return ("GTX");
      end if;
  end function;

  constant PCIE_GT_DEVICE : string := set_pcie_gt_device (C_FAMILY);

  --------------------------------------------------------------------------------
  
    function rp_interrupt_fifo_depth (C_INT_FIFO_DEPTH : integer) return integer is
    begin
      if(C_INT_FIFO_DEPTH = 0) then
        return(4);
      elsif(C_INT_FIFO_DEPTH = 1) then
        return(5);
      else
        return(6);
      end if;
  end function;

  constant PTR_WIDTH : integer  := rp_interrupt_fifo_depth (C_INT_FIFO_DEPTH);

  function family_axi_enhanced (C_FAMILY : string) return string is
    begin
      if(C_FAMILY = "virtex6") then
        return("V6");
      elsif(C_FAMILY = "spartan6") then
        return("S6");
      elsif(C_FAMILY = "7series") then
        return("X7");
      else
        return(C_FAMILY);
      end if;
  end function;

  constant FAMILY : string  := family_axi_enhanced (C_FAMILY_I);
  
  
  --------------------------------------------------------------------------------
  

  function family_user_clock (C_FAMILY, DEV, SPD : string) return integer is
    begin
      if(C_FAMILY = "virtex6") then
        return(2);
      elsif(C_FAMILY = "spartan6") then
        return(1);
      -- use DEV instead of C_FAMILY for zynq devices check
      -- clock down user_clk frequency in Zynq to help ease timing for smaller -1 devices
      -- No Gen2 support for -1 devices
      elsif(DEV = "zynq" and (SPD = "-1" or SPD = "-1i" or SPD = "-1q" or SPD = "-1l" or SPD = "-1ql" or SPD = "-1il")) then
        if (C_NO_OF_LANES = 1 or (C_NO_OF_LANES = 2 and C_MAX_LINK_SPEED = 0)) then
          if (C_S_AXI_DATA_WIDTH = 128) then
            return(2);
          else
            return (1);
          end if;
        -- This is for x2g2, x4g1/2, and x8g1/2 case which requires 125MHz at a minimum
        else
          if (C_S_AXI_DATA_WIDTH = 128) then
            return(3);
          else
            return(2);
          end if;
        end if;
      elsif (C_FAMILY = "7series") then
        if (C_S_AXI_DATA_WIDTH = 128) then
          return(3);
        elsif (C_NO_OF_LANES = 1 and C_MAX_LINK_SPEED = 0) then
          return (1);
        else
          return(2);
        end if;
      else
        return(0);
      end if;
  end function;

  --------------------------------------------------------------------------------


  function family_pcie_cap_capability_version(C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "virtex6" or C_FAMILY = "7series") then
        return(2);
      elsif(C_FAMILY = "spartan6") then
        return(1);
      else
        return(0);
      end if;
  end function;
  
  
  constant USER_CLK_FREQ : integer  := family_user_clock (C_FAMILY_I, C_FAMILY, C_SPEED);              -- 7-Series/Z(128) = 3; Z -1 half freq on x1/x2, 7-Series/V6/Z(64) = 2, S6 = 1
  constant PCIE_CAP_CAPABILITY_VERSION : integer := family_pcie_cap_capability_version (C_FAMILY_I);   -- 7-Series/V6/Z = 2, S6 = 1


  --------------------------------------------------------------------------------


  function family_total_credits_nph (C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "virtex6" or C_FAMILY = "7series") then
        return(12);
      elsif(C_FAMILY = "spartan6") then
        return(8);
      else
        return(0);
      end if;
  end function;

  constant VC0_TOTAL_CREDITS_NPH : integer := family_total_credits_nph (C_FAMILY_I);     -- V6/7-Series/Z = 12, S6 = 8

  --------------------------------------------------------------------------------
  

  function family_total_credits_pd (C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "virtex6") then
        return(154);
      elsif(C_FAMILY = "7series") then 
        return(181);        
      elsif(C_FAMILY = "spartan6") then
        return(211);
      else
        return(0);
      end if;
  end function;

  constant VC0_TOTAL_CREDITS_PD : integer := family_total_credits_pd (C_FAMILY_I);     -- V6 = 154, S6 = 211, 7-Series/Z = 181


  --------------------------------------------------------------------------------


  function family_total_credits_cd(C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "virtex6") then
        return(154);
      elsif(C_FAMILY = "7series") then 
        return(205);        
      elsif(C_FAMILY = "spartan6") then
        return(211);
      else
        return(0);
      end if;
  end function;

  constant VC0_TOTAL_CREDITS_CD : integer := family_total_credits_cd (C_FAMILY_I);     -- V6 = 154, S6 = 211, 7-Series/Z = 205


  --------------------------------------------------------------------------------


  function family_total_credits_ch(C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "virtex6" or C_FAMILY = "7series") then
        return(36);
      elsif(C_FAMILY = "spartan6") then
        return(40);
      else
        return(0);
      end if;
  end function;

  constant VC0_TOTAL_CREDITS_CH : integer := family_total_credits_ch (C_FAMILY_I);     -- V6/7-Series/Z= 36, S6 = 40


  --------------------------------------------------------------------------------


  function family_rx_ram_limit(C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "spartan6") then
        return(conv_integer(x"7ff"));
      elsif(C_FAMILY = "virtex6" or C_FAMILY = "7series") then
        return(conv_integer(x"3ff"));
      else
        return(0);
      end if;
  end function;

  constant VC0_RX_RAM_LIMIT : integer := family_rx_ram_limit (C_FAMILY_I);     -- S6 = 7FFh, V6/7-Series/Z = 3FFh


  --------------------------------------------------------------------------------


  function incl_rc_msi_cap_pvm(C_INCLUDE_RC : integer) return string is
    begin 
      if(C_INCLUDE_RC = 1) then
        return("TRUE");
      else
        return("FALSE");
      end if;
  end function;

  constant MSI_CAP_PER_VECTOR_MASKING_CAPABLE : string := incl_rc_msi_cap_pvm (C_INCLUDE_RC); -- C_INCLUDE_RC = 1 ->"TRUE" 


  --------------------------------------------------------------------------------


  function incl_rc_pcie_cap_device_port_type(C_INCLUDE_RC : integer) return integer is
    begin
      if(C_INCLUDE_RC = 1) then
        return(conv_integer(x"4"));
      else
        return(conv_integer(x"0"));
      end if;
  end function;

  constant PCIE_CAP_DEVICE_PORT_TYPE : integer := incl_rc_pcie_cap_device_port_type (C_INCLUDE_RC); --RC = 0x4, EP = 0x0


  --------------------------------------------------------------------------------

  function family_ll_replay_timeout(C_FAMILY : string) return integer is
    begin
      if (C_FAMILY = "virtex6") then
        return(conv_integer(x"0026"));
      elsif (C_FAMILY = "7series") then
        return(conv_integer(x"0000"));
      elsif (C_FAMILY = "spartan6") then
        return(conv_integer(x"00FF"));
      else
        return(0);
      end if;
  end function;

  constant LL_REPLAY_TIMEOUT : integer := family_ll_replay_timeout (C_FAMILY_I);
  
  --------------------------------------------------------------------------------


  function family_ll_replay_timeout_en (C_FAMILY : string) return string is
    begin
      if (C_FAMILY = "7series") then
        return("FALSE");
      else
        return("TRUE");
      end if;
  end function;

  constant LL_REPLAY_TIMEOUT_EN : string := family_ll_replay_timeout_en (C_FAMILY_I);     -- 7-Series/Z = "FALSE", V6/S6 = "TRUE"


  --------------------------------------------------------------------------------

  function family_pipe_pipeline_stages(C_FAMILY : string) return integer is
    begin
      if(C_FAMILY = "virtex6" or C_FAMILY = "spartan6") then
        return(0);
      elsif(C_FAMILY = "7series") then
        return(1);
      else
        return(0);
      end if;
  end function;

  constant PIPE_PIPELINE_STAGES : integer := family_pipe_pipeline_stages (C_FAMILY_I);    -- 7-Series/Z = 1, V6/S6 = 0


  --------------------------------------------------------------------------------


  function data_width_trn_dw(C_S_AXI_DATA_WIDTH : integer) return string is
    begin
      if (C_S_AXI_DATA_WIDTH = 128) then
        return("TRUE");
      else
        return("FALSE");
      end if;
  end function;

  constant TRN_DW : string := data_width_trn_dw (C_S_AXI_DATA_WIDTH);


  --------------------------------------------------------------------------------

  function data_width_user_clk2_div2(C_S_AXI_DATA_WIDTH : integer) return string is
    begin
      if(C_S_AXI_DATA_WIDTH = 128) then
        return("TRUE");
      else
        return("FALSE");
      end if;
  end function;

  constant USER_CLK2_DIV2 : string := data_width_user_clk2_div2(C_S_AXI_DATA_WIDTH);


  --------------------------------------------------------------------------------

  -- CR # 646225
  -- Move function to top level of IP
  function calc_axiread_num (C_S_AXI_DATA_WIDTH : integer) return integer is
  begin
     if C_S_AXI_DATA_WIDTH = 128 then
        return(4);
     else
        return(8);
     end if;
  end function;

  constant C_AXIREAD_NUM           : integer := calc_axiread_num (C_S_AXI_DATA_WIDTH);


  --------------------------------------------------------------------------------
  --------------------------------------------------------------------------------

  function calc_ep_link_partner_rcb (C_INCLUDE_RC, C_EP_LINK_PARTNER_RCB : integer) return integer is
  begin
     if C_INCLUDE_RC = 1 then
        return(1);
     else
        return(C_EP_LINK_PARTNER_RCB);
     end if;
  end function;

  constant EP_LINK_PARTNER_RCB     : integer := calc_ep_link_partner_rcb (C_INCLUDE_RC,C_EP_LINK_PARTNER_RCB);

-- coverage on



-- Signals

   signal axi_areset                      : std_logic;
   signal axi_aclk_in                     : std_logic;
   signal axi_ctl_aclk_in                 : std_logic;
   signal sig_axi_aclk_out                : std_logic;
   signal sig_axi_ctl_aclk_out            : std_logic;
   signal sig_pci_exp_txp                 : std_logic_vector(C_NO_OF_LANES-1 downto 0):= ZEROS(C_NO_OF_LANES-1 downto 0);
   signal sig_pci_exp_txn                 : std_logic_vector(C_NO_OF_LANES-1 downto 0):= ZEROS(C_NO_OF_LANES-1 downto 0);

   signal sig_pci_exp_rxp                 : std_logic_vector(C_NO_OF_LANES-1 downto 0);
   signal sig_pci_exp_rxn                 : std_logic_vector(C_NO_OF_LANES-1 downto 0);

   -- AXIS Write Requester Channel
   signal sig_m_axis_rw_tdata         : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
   signal sig_m_axis_rw_tstrb         : std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
   signal sig_m_axis_rw_tlast         : std_logic;
   signal sig_m_axis_rw_tvalid        : std_logic;
   signal sig_m_axis_rw_tready        : std_logic;

   -- AXIS Read Requester Channel
   signal sig_m_axis_rr_tdata         : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
   signal sig_m_axis_rr_tstrb         : std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
   signal sig_m_axis_rr_tlast         : std_logic;
   signal sig_m_axis_rr_tvalid        : std_logic;
   signal sig_m_axis_rr_tready        : std_logic;

   -- AXIS Completion Requester Channel
   signal sig_s_axis_rc_tdata         : std_logic_vector(C_M_AXIS_DATA_WIDTH-1 downto 0);
   signal sig_s_axis_rc_tstrb         : std_logic_vector(C_M_AXIS_DATA_WIDTH/8-1 downto 0);
   signal sig_s_axis_rc_tlast         : std_logic;
   signal sig_s_axis_rc_tvalid        : std_logic;
   signal sig_s_axis_rc_tready        : std_logic;

   -- AXIS Write Completer Channel
   signal sig_s_axis_cw_tdata         : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
   signal sig_s_axis_cw_tstrb         : std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
   signal sig_s_axis_cw_tlast         : std_logic;
   signal sig_s_axis_cw_tvalid        : std_logic;
   signal sig_s_axis_cw_tready        : std_logic;
   signal sig_s_axis_cw_tuser         : std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0);
      
   -- AXIS Read Completer Channel
   signal sig_s_axis_cr_tdata         : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
   signal sig_s_axis_cr_tstrb         : std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
   signal sig_s_axis_cr_tlast         : std_logic;
   signal sig_s_axis_cr_tvalid        : std_logic;
   signal sig_s_axis_cr_tready        : std_logic;
   signal sig_s_axis_cr_tuser         : std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0);

   -- AXIS Completion Completer Channel
   signal sig_m_axis_cc_tdata         : std_logic_vector(C_S_AXIS_DATA_WIDTH-1 downto 0);
   signal sig_m_axis_cc_tstrb         : std_logic_vector(C_S_AXIS_DATA_WIDTH/8-1 downto 0);
   signal sig_m_axis_cc_tlast         : std_logic;
   signal sig_m_axis_cc_tvalid        : std_logic;
   signal sig_m_axis_cc_tready        : std_logic;
   signal sig_m_axis_cc_tuser         : std_logic_vector(C_S_AXIS_USER_WIDTH-1 downto 0);

   -- AXI-Lite Slave IPIC
   signal sig_IP2Bus_Data             : std_logic_vector(31 downto 0);
   signal sig_IP2Bus_WrAck            : std_logic;
   signal sig_IP2Bus_RdAck            : std_logic;
   signal sig_IP2Bus_Error            : std_logic;
   signal sig_Bus2IP_Addr             : std_logic_vector(32-1 downto 0);
   signal sig_Bus2IP_Data             : std_logic_vector(31 downto 0);
   signal sig_Bus2IP_RNW              : std_logic;
   signal sig_Bus2IP_BE               : std_logic_vector(32/8-1 downto 0);
   signal sig_Bus2IP_CS               : std_logic;

   -- AXI-S Block Interface
   signal sig_blk_lnk_up              : std_logic;
   signal sig_blk_bus_number          : std_logic_vector(7 downto 0);
   signal sig_blk_device_number       : std_logic_vector(4 downto 0);
   signal sig_blk_function_number     : std_logic_vector(2 downto 0);
   signal sig_blk_command             : std_logic_vector(15 downto 0);
   signal sig_blk_dcontrol            : std_logic_vector(15 downto 0);
   signal sig_blk_lstatus             : std_logic_vector(15 downto 0);

   --Interrupt Strobes
   signal sig_SUR_int                 : std_logic;
   signal sig_SUC_int                 : std_logic;
   signal sig_SCT_int                 : std_logic;
   signal sig_SEP_int                 : std_logic;
   signal sig_SCA_int                 : std_logic;
   signal sig_SIB_int                 : std_logic;
   signal sig_MDE_int                 : std_logic;
   signal sig_MSE_int                 : std_logic;
   signal sig_MEP_int                 : std_logic;
   --signal sig_MLE_int                 : std_logic;
   --signal sig_MEC_int                 : std_logic;
   signal interrupt_vector            : std_logic_vector(NUM_OF_INTERRUPTS-1 downto 0);
   signal np_cpl_pending              : std_logic;
   signal np_cpl_pending_qual         : std_logic;
   signal sig_blk_interrupt           : std_logic;
   signal sig_blk_interrupt_rdy       : std_logic;
   signal sig_blk_interrupt_assert    : std_logic;
   signal sig_blk_interrupt_di        : std_logic_vector(7 downto 0);
   signal sig_blk_interrupt_msienable : std_logic;
   signal sig_intx_msi_request        : std_logic;
   signal sig_intx_msi_grant          : std_logic;
   signal sig_msi_vector_num          : std_logic_vector(4 downto 0);
   signal intx_msi_request_1d         : std_logic;
   signal intx_msi_request_2d         : std_logic;
   signal intx_msi_request_3d         : std_logic;
   signal msi_vector_num_1d           : std_logic_vector(4 downto 0);
   signal msi_vector_num_2d           : std_logic_vector(4 downto 0);
   signal sig_mmcm_lock               : std_logic;
   signal RP_bridge_en                : std_logic;

   type legint_msiSM_STATES is (NO_INTR,
                                INTR_HS);
   signal legint_msiSM : legint_msiSM_STATES;
   signal INTX_state                  : std_logic;
   constant SELECTED_INT              : std_logic_vector(7 downto 0) := conv_std_logic_vector(C_INTERRUPT_PIN-1, 8);

   signal counter_50: integer := 0;

-- Signals for np_req_mode: if C_TRN_NP_FC = "TRUE"
   signal sig_rx_np_req               : std_logic;
   signal rx_np_req_cntr              : integer range 0 to 15;
   signal np_pkt_complete             : std_logic_vector(1 downto 0); -- bit[1] = rdndreqpipeline; bit[0] = rdreqpipeline
-- End np_req_mode signals

-- Signals for np_ok_mode: if C_TRN_NP_FC = "FALSE"
   type rx_np_okSM_STATES is (INIT,
                              WAIT_PIPE_LATENCY,
                              CHECK_NP_PIPELINE,
                              ASSERT_NP_OK);
   signal rx_np_okSM                  : rx_np_okSM_STATES;
   constant RX_PIPE_LATENCY           : integer := 12;
   signal sig_rx_np_ok                : std_logic;
   signal rx_np_ok_int                : std_logic;
   signal rx_np_ok_cntr               : integer range 0 to 15;
   signal pipe_latency_cntr           : integer range 0 to 15;
   signal disable_rx_np_ok            : std_logic;
   signal rdndreqpipeline             : std_logic_vector(2 downto 0);
   signal rdreqpipeline               : std_logic_vector(2 downto 0);
   signal rdndreqpipeline_d           : std_logic_vector(2 downto 0);
   signal rdreqpipeline_d             : std_logic_vector(2 downto 0);
-- End np_ok_mode signals

   signal config_gen_req              : std_logic;

begin

   -- Tx
   pci_exp_txp                   <= sig_pci_exp_txp;
   pci_exp_txn                   <= sig_pci_exp_txn;
   -- Rx
   sig_pci_exp_rxp               <= pci_exp_rxp;
   sig_pci_exp_rxn               <= pci_exp_rxn;
   
   axi_areset                    <= not(axi_aresetn);
clk_input : if AXI_ACLK_LOOPBACK = "TRUE" generate
   axi_aclk_in			 <= axi_aclk;
   axi_ctl_aclk_in               <= axi_ctl_aclk;
end generate;
intrnl_clk_input : if AXI_ACLK_LOOPBACK = "FALSE" generate
   axi_aclk_in			 <= sig_axi_aclk_out;
   axi_ctl_aclk_in               <= sig_axi_ctl_aclk_out;
end generate;
   axi_aclk_out			 <= sig_axi_aclk_out;
   axi_ctl_aclk_out              <= sig_axi_ctl_aclk_out;

   interrupt_vector              <= sig_MEP_int & sig_MSE_int & sig_MDE_int & sig_SIB_int & sig_SCA_int & sig_SEP_int & sig_SCT_int & sig_SUC_int & sig_SUR_int;
   MSI_enable                    <= sig_blk_interrupt_msienable;
   INTX_MSI_Grant                <= sig_intx_msi_grant;
   sig_intx_msi_request          <= INTX_MSI_Request;
   sig_msi_vector_num            <= MSI_Vector_Num;
   np_cpl_pending_qual           <= np_cpl_pending when C_INCLUDE_RC = 1 else '1';

   mmcm_lock                     <= sig_mmcm_lock;
   user_link_up                  <= sig_blk_lnk_up;

np_req_mode: if C_TRN_NP_FC = "TRUE" generate begin
   sig_rx_np_ok            <= '0';

--**************************************************************************************************
-- This StateMachine will actively look for available NP Buffer space of MM/S MasterBridge Rd module
-- and make full use of rx_np_req signal to control NP traffic on receive side. Hence avoids potential
-- PCIe-Rx MemRd buffer overflow problem
--**************************************************************************************************

   rx_np_req_proc : process (axi_aclk_in)
   begin
      if(rising_edge(axi_aclk_in)) then
         if(axi_aresetn = '0' or sig_blk_lnk_up = '0') then
            sig_rx_np_req            <= '0';
            
            -- 128-bit: assert rx_np_req for 4 clock cycles, doing so will accept up to 4 NP packets
            -- if it has any
            if C_S_AXI_DATA_WIDTH = 128 then -- 128-bit
                rx_np_req_cntr   <= 4;

            -- 64-bit: assert rx_np_req for 5 clock cycles, doing so will accept up to 5 NP packets
            -- if it has any
            elsif C_S_AXI_DATA_WIDTH = 64 then -- 64-bit
                rx_np_req_cntr   <= 5;

            -- 32-bit: assert rx_np_req for 9 clock cycles, doing so will accept up to 9 NP packets
            -- if it has any
            else -- 32-bit
                rx_np_req_cntr   <= 9;
            end if; -- C_S_AXI_DATA_WIDTH
            
         else
            
            -- Request more NP packet if the pipeline still have some space
            if rx_np_req_cntr /= 0 then
                sig_rx_np_req    <= '1';
            else
                sig_rx_np_req    <= '0';
            end if;
            
            if np_pkt_complete(0) = '1' or np_pkt_complete(1) = '1' then
	        -- OR'ing because it can only be completion with data or without data but not both
                -- Increment one when completion is sent (a read request has been serviced), and
                --  there's no pending rx_np_req signal update
                -- If there's pending update, then it will be +1 then -1, so no change
                if rx_np_req_cntr = 0 then
                    rx_np_req_cntr   <= rx_np_req_cntr + 1;
                end if;
            else
                -- Decrement one if there's pending update
                if rx_np_req_cntr /= 0 then
                    rx_np_req_cntr   <= rx_np_req_cntr - 1;
                end if;
            end if;
            
         end if; -- axi_areset
      end if; -- axi_aclk
   end process;
end generate;

np_ok_mode: if C_TRN_NP_FC = "FALSE" generate begin
   disable_rx_np_ok              <= '1' when rdreqpipeline_d = "000" and rdndreqpipeline_d = "000" and sig_s_axis_cr_tlast = '1' else '0';
   sig_rx_np_ok                  <= rx_np_ok_int and (not(disable_rx_np_ok)) when C_S_AXI_DATA_WIDTH = 128 else rx_np_ok_int;
   sig_rx_np_req                 <= '1';

--**************************************************************************************************
-- This StateMachine will actively look for available NP Buffer space of MM/S MasterBridge Rd module
-- and make full use of rx_np_ok signal to control NP traffic on receive side. Hence avoids potential
-- PCIe-Rx Cpl buffer overflow problem
--**************************************************************************************************

   rx_np_ok_proc : process (axi_aclk_in)
   begin
      if(rising_edge(axi_aclk_in)) then
         if(axi_aresetn = '0') then
            rx_np_ok_int              <= '0';
            rx_np_ok_cntr             <= 0;
            pipe_latency_cntr         <= 0;
            rdreqpipeline_d           <= "000";
            rdndreqpipeline_d         <= "000";
            rx_np_okSM                <= INIT;
         else
            rdreqpipeline_d           <= rdreqpipeline;
            rdndreqpipeline_d         <= rdndreqpipeline;
            
            case rx_np_okSM is
            
            when INIT =>

               rx_np_ok_cntr      <= rx_np_ok_cntr;
	       pipe_latency_cntr  <= pipe_latency_cntr;
               -- De-assert rx_np_ok as soon as 1st NP TLP on CR interface is encountered
               -- Assumption here is pessimistic becuase there can be many back-2-back MRds
               -- In 128-bit mode, situation is worse as there could be 5 MRd back-to-back
               -- even if we de-assert rx_np_ok after encountering 1st NP TLP on CR interface
               if rdreqpipeline_d = "000" and rdndreqpipeline_d = "000" and 
                  sig_s_axis_cr_tlast = '1' then
                  rx_np_ok_int     <= '0';
                  rx_np_okSM       <= WAIT_PIPE_LATENCY;
               else
                  rx_np_ok_int     <= '1';
               end if;

            -- Wait for enough amout of time so that NP TLPs can propagate from Block to MM/S masterbridge rd
            -- and rdreqpipeline gets updated
            when WAIT_PIPE_LATENCY =>

               rx_np_ok_cntr        <= rx_np_ok_cntr;
               rx_np_ok_int         <= rx_np_ok_int;
               -- RX_PIPE_LATENCY is constant which is set to 12 based on best practices and assumption
               -- that MRds in-flight along with those block may give even after de-asserting rx_np_ok will be
               -- pipelined in MM/S masterbridge rd module successfully
               if pipe_latency_cntr = RX_PIPE_LATENCY then
                  rx_np_okSM        <= CHECK_NP_PIPELINE;
                  pipe_latency_cntr <= 0;
               else
                  pipe_latency_cntr <= pipe_latency_cntr + 1;
               end if;

            -- Check if there is some slot vacant to accomodate more MRd
            when CHECK_NP_PIPELINE =>

               pipe_latency_cntr   <= pipe_latency_cntr;
	       -- Pipeline is found empty... go to INIT state
               if rdreqpipeline_d = "000" and rdndreqpipeline_d = "000" then
                  rx_np_okSM       <= INIT;
                  rx_np_ok_int     <= '1';

               -- Pipeline is not empty but can accomodate more TLPs
               -- At this point, MM/S masterbridge rd can accomodate 3 additional NP TLP in 32/64-bit mode
               -- and 4 NP TLPs in 128-bit mode
               elsif rdreqpipeline_d = "001" or rdndreqpipeline_d = "001" then

                  -- 128-bit: assert rx_np_ok for 4 clock cycles and by doing so, block may throw 4 NP TLPs
                  -- if it will have any
                  if C_S_AXI_DATA_WIDTH = 128 then -- 128-bit
                     rx_np_ok_cntr    <= 4;

                  -- 64-bit: assert rx_np_ok for 6 clock cycles and by doing so, block may throw 3 NP TLPs
                  -- if it will have any
                  elsif C_S_AXI_DATA_WIDTH = 64 then -- 64-bit
                     rx_np_ok_cntr    <= 6;

                  -- 32-bit: assert rx_np_ok for 9 clock cycles and by doing so, block may throw 3 NP TLPs
                  -- if it will have any
                  else -- 32-bit
                     rx_np_ok_cntr    <= 9;
                  end if;

                  rx_np_okSM       <= ASSERT_NP_OK;

               -- At this point, MM/S masterbridge rd can accomodate 2 additional NP TLP in 32/64-bit mode
               -- and 3 NP TLPs in 128-bit mode
               elsif rdreqpipeline_d = "010" or rdndreqpipeline_d = "010" then

                  -- 32-bit: assert rx_np_ok for 6 clock cycles and by doing so, block may throw 2 NP TLPs
                  -- if it will have any
                  if C_S_AXI_DATA_WIDTH = 32 then -- 32-bit
                     rx_np_ok_cntr    <= 6;

                  -- 64/128-bit: assert rx_np_ok for 3 clock cycles and by doing so, block may throw 
                  -- 3 NP TLPs in 128-bit mode and 2 TLPs in 64-bit mode if it will have any
                  else -- 64/128-bit
                     rx_np_ok_cntr    <= 3;
                  end if;

                  rx_np_okSM       <= ASSERT_NP_OK;

               -- At this point, MM/S masterbridge rd can accomodate 1 additional NP TLP in 32/64-bit mode
               -- and 2 NP TLPs in 128-bit mode
               elsif rdreqpipeline_d = "011" or rdndreqpipeline_d = "011" then
                  rx_np_okSM       <= ASSERT_NP_OK;
                  rx_np_ok_cntr    <= 2;
               end if;

            -- SM will come to this state when rdreqpipeline will have available space sufficient enough to
            -- accomodate 1 or more MRd TLPs. This state retains rx_np_ok asserted for number of clock cycles
            -- programmed in rx_np_ok_cntr before next check iteration
            when ASSERT_NP_OK =>

               pipe_latency_cntr   <= pipe_latency_cntr;
	       if rx_np_ok_cntr = 0 then
                  rx_np_okSM       <= WAIT_PIPE_LATENCY;
                  rx_np_ok_int     <= '0';
               else
                  rx_np_ok_cntr    <= rx_np_ok_cntr - 1;
                  rx_np_ok_int     <= '1';
               end if;

            end case;

         end if;
      end if;
   end process;
end generate;

--***************************************************************************************************
-- Legacy and MSI interrupt logic
--***************************************************************************************************

   legacy_MSI_interrupt_proc : process (axi_aclk_in)
   begin
      if(rising_edge(axi_aclk_in)) then
         if(axi_aresetn = '0') then
            sig_blk_interrupt         <= '0';
            sig_blk_interrupt_assert  <= '0';
            sig_blk_interrupt_di      <= (others => '0');
            INTX_state                <= '0';
            legint_msiSM              <= NO_INTR;
            intx_msi_request_1d       <= '0';
            intx_msi_request_2d       <= '0';
            intx_msi_request_3d       <= '0';
            msi_vector_num_1d         <= (others => '0');
            msi_vector_num_2d         <= (others => '0');
            sig_intx_msi_grant        <= '0';
         elsif C_INCLUDE_RC = 0 then -- only for End Point
            intx_msi_request_1d       <= sig_intx_msi_request;
            intx_msi_request_2d       <= intx_msi_request_1d;
            intx_msi_request_3d       <= intx_msi_request_2d;
            msi_vector_num_1d         <= sig_msi_vector_num;
            msi_vector_num_2d         <= msi_vector_num_1d;
            case legint_msiSM is

               when NO_INTR =>
                  if sig_blk_interrupt_msienable = '1' then
                     if intx_msi_request_2d = '1' and intx_msi_request_3d = '0' then --positive edge detect
                        sig_blk_interrupt         <= '1';
                        sig_blk_interrupt_assert  <= '0';
                        sig_blk_interrupt_di      <= ("000" & msi_vector_num_2d);
                        legint_msiSM              <= INTR_HS;
                     end if;
                  else
                     if sig_intx_msi_request /= INTX_state then
                        sig_blk_interrupt         <= '1';
                        sig_blk_interrupt_assert  <= sig_intx_msi_request;
                        sig_blk_interrupt_di      <= SELECTED_INT;
                        INTX_state                <= sig_intx_msi_request;
                        legint_msiSM              <= INTR_HS;
                     end if;
                  end if;
                  sig_intx_msi_grant  <= '0';

               when INTR_HS =>
                  INTX_state                   <= INTX_state;
		  if sig_blk_interrupt_rdy = '1' then
                     sig_blk_interrupt         <= '0';
                     sig_blk_interrupt_assert  <= '0';
                     sig_blk_interrupt_di      <= (others => '0');
                     legint_msiSM              <= NO_INTR;
                     sig_intx_msi_grant        <= '1';
                  end if;

            end case;
         end if;
      end if;
   end process;

   comp_axi_pcie_mm_s: entity axi_pcie_v2_9_14.axi_pcie_mm_s
    generic map(
      --Family Generics
      -- C_FAMILY                      => C_FAMILY_I,
      C_FAMILY                      => C_FAMILY,  -- MM/S bridge gets derivative C_FAMILY parameter      
      C_S_AXI_ID_WIDTH              => C_S_AXI_ID_WIDTH,
      --C_M_AXI_THREAD_ID_WIDTH       => C_M_AXI_THREAD_ID_WIDTH,
      C_S_AXI_ADDR_WIDTH            => C_S_AXI_ADDR_WIDTH,
      C_S_AXI_DATA_WIDTH            => C_S_AXI_DATA_WIDTH,
      C_M_AXI_ADDR_WIDTH            => C_M_AXI_ADDR_WIDTH,
      C_M_AXI_DATA_WIDTH            => C_M_AXI_DATA_WIDTH,
      C_S_AXIS_DATA_WIDTH           => C_S_AXIS_DATA_WIDTH,
      C_M_AXIS_DATA_WIDTH           => C_M_AXIS_DATA_WIDTH,
      C_COMP_TIMEOUT                => C_COMP_TIMEOUT,
      C_USER_CLK_FREQ               => USER_CLK_FREQ,
      C_USER_CLK2_DIV2              => USER_CLK2_DIV2,
      C_INCLUDE_RC                  => C_INCLUDE_RC,
      C_S_AXI_SUPPORTS_NARROW_BURST => C_S_AXI_SUPPORTS_NARROW_BURST,
      C_EP_LINK_PARTNER_RCB         => EP_LINK_PARTNER_RCB,
      C_INCLUDE_BAROFFSET_REG       => C_INCLUDE_BAROFFSET_REG,
      C_AXIREAD_NUM                 => C_AXIREAD_NUM,   -- CR # 646225
      C_AXIBAR_NUM                  => C_AXIBAR_NUM,
      C_AXIBAR2PCIEBAR_0            => C_AXIBAR2PCIEBAR_0,
      C_AXIBAR2PCIEBAR_1            => C_AXIBAR2PCIEBAR_1,
      C_AXIBAR2PCIEBAR_2            => C_AXIBAR2PCIEBAR_2,
      C_AXIBAR2PCIEBAR_3            => C_AXIBAR2PCIEBAR_3,
      C_AXIBAR2PCIEBAR_4            => C_AXIBAR2PCIEBAR_4,
      C_AXIBAR2PCIEBAR_5            => C_AXIBAR2PCIEBAR_5,
      C_AXIBAR_AS_0                 => C_AXIBAR_AS_0,
      C_AXIBAR_AS_1                 => C_AXIBAR_AS_1,
      C_AXIBAR_AS_2                 => C_AXIBAR_AS_2,
      C_AXIBAR_AS_3                 => C_AXIBAR_AS_3,
      C_AXIBAR_AS_4                 => C_AXIBAR_AS_4,
      C_AXIBAR_AS_5                 => C_AXIBAR_AS_5,
      C_AXIBAR_0                    => C_AXIBAR_0,
      C_AXIBAR_HIGHADDR_0           => C_AXIBAR_HIGHADDR_0,
      C_AXIBAR_1                    => C_AXIBAR_1,
      C_AXIBAR_HIGHADDR_1           => C_AXIBAR_HIGHADDR_1,
      C_AXIBAR_2                    => C_AXIBAR_2,
      C_AXIBAR_HIGHADDR_2           => C_AXIBAR_HIGHADDR_2,
      C_AXIBAR_3                    => C_AXIBAR_3,
      C_AXIBAR_HIGHADDR_3           => C_AXIBAR_HIGHADDR_3,
      C_AXIBAR_4                    => C_AXIBAR_4,
      C_AXIBAR_HIGHADDR_4           => C_AXIBAR_HIGHADDR_4,
      C_AXIBAR_5                    => C_AXIBAR_5,
      C_AXIBAR_HIGHADDR_5           => C_AXIBAR_HIGHADDR_5,
      C_PCIEBAR_NUM                 => C_PCIEBAR_NUM,
      C_PCIEBAR_AS                  => C_PCIEBAR_AS,
      C_PCIEBAR_LEN_0               => C_PCIEBAR_LEN_0,
      C_PCIEBAR2AXIBAR_0            => C_PCIEBAR2AXIBAR_0,
      C_PCIEBAR2AXIBAR_0_SEC        => C_PCIEBAR2AXIBAR_0_SEC,
      C_PCIEBAR_LEN_1               => C_PCIEBAR_LEN_1,
      C_PCIEBAR2AXIBAR_1            => C_PCIEBAR2AXIBAR_1,
      C_PCIEBAR2AXIBAR_1_SEC        => C_PCIEBAR2AXIBAR_1_SEC,
      C_PCIEBAR_LEN_2               => C_PCIEBAR_LEN_2,
      C_PCIEBAR2AXIBAR_2            => C_PCIEBAR2AXIBAR_2,
      C_PCIEBAR2AXIBAR_2_SEC        => C_PCIEBAR2AXIBAR_2_SEC,
      C_S_AXIS_USER_WIDTH           => C_S_AXIS_USER_WIDTH,
      C_TRN_NP_FC                   => C_TRN_NP_FC,
      C_AXIBAR_CHK_SLV_ERR          => C_AXIBAR_CHK_SLV_ERR
    )
    port map(
      -- AXI Global
      axi_aclk                => axi_aclk_in,
      reset                   => axi_aresetn,

      -- AXI Slave Write Address Channel
      s_axi_awid              => s_axi_awid,
      s_axi_awaddr            => s_axi_awaddr,
      s_axi_awregion          => s_axi_awregion,
      s_axi_awlen             => s_axi_awlen,
      s_axi_awsize            => s_axi_awsize,
      s_axi_awburst           => s_axi_awburst,
      s_axi_awvalid           => s_axi_awvalid,
      s_axi_awready           => s_axi_awready,

      -- AXI Slave Write Data Channel
      s_axi_wdata             => s_axi_wdata,
      s_axi_wstrb             => s_axi_wstrb,
      s_axi_wlast             => s_axi_wlast,
      s_axi_wvalid            => s_axi_wvalid,
      s_axi_wready            => s_axi_wready,

      -- AXI Slave Write Response Channel
      s_axi_bid               => s_axi_bid,
      s_axi_bresp             => s_axi_bresp,
      s_axi_bvalid            => s_axi_bvalid,
      s_axi_bready            => s_axi_bready,

      -- AXI Slave Read Address Channel
      s_axi_arid              => s_axi_arid,
      s_axi_araddr            => s_axi_araddr,
      s_axi_arregion          => s_axi_arregion,
      s_axi_arlen             => s_axi_arlen,
      s_axi_arsize            => s_axi_arsize,
      s_axi_arburst           => s_axi_arburst,
      s_axi_arvalid           => s_axi_arvalid,
      s_axi_arready           => s_axi_arready,

      -- AXI Slave Read Data Channel
      s_axi_rid               => s_axi_rid,
      s_axi_rdata             => s_axi_rdata,
      s_axi_rresp             => s_axi_rresp,
      s_axi_rlast             => s_axi_rlast,
      s_axi_rvalid            => s_axi_rvalid,
      s_axi_rready            => s_axi_rready,

      -- AXIS Write Requester Channel
      m_axis_rw_tdata         => sig_m_axis_rw_tdata,
      m_axis_rw_tstrb         => sig_m_axis_rw_tstrb,
      m_axis_rw_tlast         => sig_m_axis_rw_tlast,
      m_axis_rw_tvalid        => sig_m_axis_rw_tvalid,
      m_axis_rw_tready        => sig_m_axis_rw_tready,

      -- AXIS Read Requester Channel
      m_axis_rr_tdata         => sig_m_axis_rr_tdata,
      m_axis_rr_tstrb         => sig_m_axis_rr_tstrb,
      m_axis_rr_tlast         => sig_m_axis_rr_tlast,
      m_axis_rr_tvalid        => sig_m_axis_rr_tvalid,
      m_axis_rr_tready        => sig_m_axis_rr_tready,

      -- AXIS Completion Requester Channel
      s_axis_rc_tdata         => sig_s_axis_rc_tdata,
      s_axis_rc_tstrb         => sig_s_axis_rc_tstrb,
      s_axis_rc_tlast         => sig_s_axis_rc_tlast,
      s_axis_rc_tvalid        => sig_s_axis_rc_tvalid,
      s_axis_rc_tready        => sig_s_axis_rc_tready,

      -- AXI Master Write Address Channel
      m_axi_awaddr            => m_axi_awaddr,
      m_axi_awlen             => m_axi_awlen,
      m_axi_awsize            => m_axi_awsize,
      m_axi_awburst           => m_axi_awburst,
      m_axi_awprot            => m_axi_awprot,
      m_axi_awvalid           => m_axi_awvalid,
      m_axi_awready           => m_axi_awready,
      --m_axi_awid              => m_axi_awid,
      m_axi_awlock            => m_axi_awlock,
      m_axi_awcache           => m_axi_awcache,

      -- AXI Master Write Data Channel
      m_axi_wdata             => m_axi_wdata,
      m_axi_wstrb             => m_axi_wstrb,
      m_axi_wlast             => m_axi_wlast,
      m_axi_wvalid            => m_axi_wvalid,
      m_axi_wready            => m_axi_wready,

      -- AXI Master Write Response Channel
      m_axi_bresp             => m_axi_bresp,
      m_axi_bvalid            => m_axi_bvalid,
      m_axi_bready            => m_axi_bready,

      -- AXI Master Read Address Channel
      --m_axi_arid              => m_axi_arid,
      m_axi_araddr            => m_axi_araddr,
      m_axi_arlen             => m_axi_arlen,
      m_axi_arsize            => m_axi_arsize,
      m_axi_arburst           => m_axi_arburst,
      m_axi_arprot            => m_axi_arprot,
      m_axi_arvalid           => m_axi_arvalid,
      m_axi_arready           => m_axi_arready,
      m_axi_arlock            => m_axi_arlock,
      m_axi_arcache           => m_axi_arcache,

      -- AXI Master Read Data Channel
      m_axi_rdata             => m_axi_rdata,
      m_axi_rresp             => m_axi_rresp,
      m_axi_rlast             => m_axi_rlast,
      m_axi_rvalid            => m_axi_rvalid,
      m_axi_rready            => m_axi_rready,

      -- AXIS Write Completer Channel
      s_axis_cw_tdata         => sig_s_axis_cw_tdata,
      s_axis_cw_tstrb         => sig_s_axis_cw_tstrb,
      s_axis_cw_tlast         => sig_s_axis_cw_tlast,
      s_axis_cw_tvalid        => sig_s_axis_cw_tvalid,
      s_axis_cw_tready        => sig_s_axis_cw_tready,
      s_axis_cw_tuser         => sig_s_axis_cw_tuser,
      
      -- AXIS Read Completer Channel
      s_axis_cr_tdata         => sig_s_axis_cr_tdata,
      s_axis_cr_tstrb         => sig_s_axis_cr_tstrb,
      s_axis_cr_tlast         => sig_s_axis_cr_tlast,
      s_axis_cr_tvalid        => sig_s_axis_cr_tvalid,
      s_axis_cr_tready        => sig_s_axis_cr_tready,
      s_axis_cr_tuser         => sig_s_axis_cr_tuser,

      -- AXIS Completion Completer Channel
      m_axis_cc_tdata         => sig_m_axis_cc_tdata,
      m_axis_cc_tstrb         => sig_m_axis_cc_tstrb,
      m_axis_cc_tlast         => sig_m_axis_cc_tlast,
      m_axis_cc_tvalid        => sig_m_axis_cc_tvalid,
      m_axis_cc_tready        => sig_m_axis_cc_tready,
      m_axis_cc_tuser         => sig_m_axis_cc_tuser,

      -- AXI-Lite Slave IPIC
      IP2Bus_Data             => sig_IP2Bus_Data,
      IP2Bus_WrAck            => sig_IP2Bus_WrAck,
      IP2Bus_RdAck            => sig_IP2Bus_RdAck,
      IP2Bus_Error            => sig_IP2Bus_Error,
      Bus2IP_Addr             => sig_Bus2IP_Addr,
      Bus2IP_Data             => sig_Bus2IP_Data,
      Bus2IP_RNW              => sig_Bus2IP_RNW,
      Bus2IP_BE               => sig_Bus2IP_BE,
      Bus2IP_CS               => sig_Bus2IP_CS,

      -- AXI-S Block Interface
      blk_lnk_up              => sig_blk_lnk_up,
      blk_bus_number          => sig_blk_bus_number,
      blk_device_number       => sig_blk_device_number,
      blk_function_number     => sig_blk_function_number,
      blk_command             => sig_blk_command,
      blk_dcontrol            => sig_blk_dcontrol,
      blk_lstatus             => sig_blk_lstatus,
      np_cpl_pending          => np_cpl_pending,-- out  std_logic;
      RP_bridge_en            => RP_bridge_en,

      --Interrupt Strobes
      SUR_int                 => sig_SUR_int,
      SUC_int                 => sig_SUC_int,
      SCT_int                 => sig_SCT_int,
      SEP_int                 => sig_SEP_int,
      SCA_int                 => sig_SCA_int,
      SIB_int                 => sig_SIB_int,
      MDE_int                 => sig_MDE_int, -- Master DECERR interrupt
      MSE_int                 => sig_MSE_int, -- Master SLVERR interrupt
      MEP_int                 => sig_MEP_int, -- Slave Error Poison interrupt
      --MLE_int                 => sig_MLE_int, -- Link Down interrupt
      --MEC_int                 => sig_MEC_int  -- ECRC Error interrupt
      
      -- signals used to keep track NP buffer availability
-- Signals for np_req_mode: if C_TRN_NP_FC = "TRUE"
      np_pkt_complete         => np_pkt_complete,
-- End np_req_mode signals
      
-- Signals for np_ok_mode: if C_TRN_NP_FC = "FALSE"
      rdndreqpipeline         => rdndreqpipeline,
      rdreqpipeline           => rdreqpipeline,
-- End np_ok_mode signals

      config_gen_req          => config_gen_req
    );

   comp_axi_enhanced_pcie: entity axi_pcie_v2_9_14.axi_enhanced_pcie
    generic map(
      C_DATA_WIDTH                             => C_S_AXIS_DATA_WIDTH,
      STRB_WIDTH                               => C_S_AXIS_DATA_WIDTH/8,
      NO_SLV_ERR                               => NO_SLV_ERR,
      BAR0_U                                   => BAR0_U,
      BAR0_L                                   => BAR0_L,
      BAR1_U                                   => BAR1_U,
      BAR1_L                                   => BAR1_L,
      BAR2_U                                   => BAR2_U,
      BAR2_L                                   => BAR2_L,
      BAR3_U                                   => BAR3_U,
      BAR3_L                                   => BAR3_L,
      BAR4_U                                   => BAR4_U,
      BAR4_L                                   => BAR4_L,
      BAR5_U                                   => BAR5_U,
      BAR5_L                                   => BAR5_L,
      CARDBUS_CIS_POINTER                      => conv_integer(x"00000000"),
      CLASS_CODE                               => conv_integer(C_CLASS_CODE),
      CMD_INTX_IMPLEMENTED                     => "TRUE",
      CPL_TIMEOUT_DISABLE_SUPPORTED            => "FALSE",
      CPL_TIMEOUT_RANGES_SUPPORTED             => conv_integer(x"0"),-- 2
      DEV_CAP_EXT_TAG_SUPPORTED                => "TRUE",
      DEV_CAP_MAX_PAYLOAD_SUPPORTED            => 1,-- 256 bytes
      DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT        => 1,
      DEVICE_ID                                => conv_integer(C_DEVICE_ID),
      DISABLE_LANE_REVERSAL                    => "TRUE",    -- CR # 618714 "FALSE",
      DISABLE_SCRAMBLING                       => "FALSE",
      DSN_BASE_PTR                             => conv_integer(x"100"),
      DSN_CAP_NEXTPTR                          => conv_integer(x"000"),
      DSN_CAP_ON                               => "TRUE",
      ENABLE_MSG_ROUTE                         => conv_integer(x"27f"),
      ENABLE_RX_TD_ECRC_TRIM                   => "TRUE",
      EXPANSION_ROM_U                          => 0,
      EXPANSION_ROM_L                          => 0, 
      EXT_CFG_CAP_PTR                          => conv_integer(x"3f"),
      EXT_CFG_XP_CAP_PTR                       => conv_integer(x"3ff"),
      HEADER_TYPE                              => C_INCLUDE_RC,
      INTERRUPT_PIN                            => C_INTERRUPT_PIN, --: integer:= conv_integer(x"00"),
      LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP   => LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP_LOCAL,
      LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP => "FALSE",
      LINK_CAP_MAX_LINK_SPEED                  => C_MAX_LINK_SPEED+1, -- 2.5 GT/s, 5.0 GT/s
      LINK_CAP_MAX_LINK_WIDTH                  => C_NO_OF_LANES,
      LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE     => "FALSE",
      LINK_CONTROL_RCB                         => 0,
      LINK_CTRL2_DEEMPHASIS                    => "FALSE",
      LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE   => "FALSE",
      LINK_CTRL2_TARGET_LINK_SPEED             => C_MAX_LINK_SPEED+1, -- 2.5 GT/s, 5.0 GT/s
      LINK_STATUS_SLOT_CLOCK_CONFIG            => C_SLOT_CLOCK_CONFIG,
      LL_ACK_TIMEOUT                           => conv_integer(x"0000"),
      LL_ACK_TIMEOUT_EN                        => "FALSE",
      LL_ACK_TIMEOUT_FUNC                      => 0,
      LL_REPLAY_TIMEOUT                        => LL_REPLAY_TIMEOUT,
      LL_REPLAY_TIMEOUT_EN                     => LL_REPLAY_TIMEOUT_EN,
      LL_REPLAY_TIMEOUT_FUNC                   => 1,
      LTSSM_MAX_LINK_WIDTH                     => C_NO_OF_LANES,
      MSI_DECODE_ENABLE                        => C_MSI_DECODE_ENABLE,
      MSI_CAP_MULTIMSGCAP                      => C_NUM_MSI_REQ,
      MSI_CAP_MULTIMSG_EXTENSION               => 0,
      MSI_CAP_ON                               => "TRUE",
      MSI_CAP_PER_VECTOR_MASKING_CAPABLE       => MSI_CAP_PER_VECTOR_MASKING_CAPABLE,
      MSI_CAP_64_BIT_ADDR_CAPABLE              => "TRUE",

      MSIX_CAP_ON                              => "FALSE",
      MSIX_CAP_PBA_BIR                         => 0,
      MSIX_CAP_PBA_OFFSET                      => conv_integer(x"00000050"),
      MSIX_CAP_TABLE_BIR                       => 0,
      MSIX_CAP_TABLE_OFFSET                    => conv_integer(x"00000040"),
      MSIX_CAP_TABLE_SIZE                      => conv_integer(x"000"),

      PCIE_CAP_DEVICE_PORT_TYPE                => PCIE_CAP_DEVICE_PORT_TYPE,
      PCIE_CAP_INT_MSG_NUM                     => conv_integer(x"00"),
      PCIE_CAP_NEXTPTR                         => conv_integer(x"00"),
      PCIE_DRP_ENABLE                          => "FALSE",
      PIPE_PIPELINE_STAGES                     => PIPE_PIPELINE_STAGES,  -- 0 - 0 stages, 1 - 1 stage, 2 - 2 stages

      PM_CAP_DSI                               => "TRUE",
      PM_CAP_D1SUPPORT                         => "FALSE",
      PM_CAP_D2SUPPORT                         => "FALSE",
      PM_CAP_NEXTPTR                           => conv_integer(x"48"),
      PM_CAP_PMESUPPORT                        => conv_integer(x"00"),
      PM_CSR_NOSOFTRST                         => "TRUE",

      PM_DATA_SCALE0                           => conv_integer(x"0"),
      PM_DATA_SCALE1                           => conv_integer(x"0"),
      PM_DATA_SCALE2                           => conv_integer(x"0"),
      PM_DATA_SCALE3                           => conv_integer(x"0"),
      PM_DATA_SCALE4                           => conv_integer(x"0"),
      PM_DATA_SCALE5                           => conv_integer(x"0"),
      PM_DATA_SCALE6                           => conv_integer(x"0"),
      PM_DATA_SCALE7                           => conv_integer(x"0"),

      PM_DATA0                                 => conv_integer(x"00"),
      PM_DATA1                                 => conv_integer(x"00"),
      PM_DATA2                                 => conv_integer(x"00"),
      PM_DATA3                                 => conv_integer(x"00"),
      PM_DATA4                                 => conv_integer(x"00"),
      PM_DATA5                                 => conv_integer(x"00"),
      PM_DATA6                                 => conv_integer(x"00"),
      PM_DATA7                                 => conv_integer(x"00"),
      REF_CLK_FREQ                             => C_REF_CLK_FREQ,-- 0 - 100 MHz, 1 - 125 MHz, 2 - 250 MHz
      REVISION_ID                              => conv_integer(C_REV_ID),
      ROOT_CAP_CRS_SW_VISIBILITY               => "FALSE",
      SPARE_BIT0                               => 0,
      SUBSYSTEM_ID                             => conv_integer(C_SUBSYSTEM_ID),
      SUBSYSTEM_VENDOR_ID                      => conv_integer(C_SUBSYSTEM_VENDOR_ID),
      SLOT_CAP_ATT_BUTTON_PRESENT              => "FALSE",
      SLOT_CAP_ATT_INDICATOR_PRESENT           => "FALSE",
      SLOT_CAP_ELEC_INTERLOCK_PRESENT          => "FALSE",
      SLOT_CAP_HOTPLUG_CAPABLE                 => "FALSE",
      SLOT_CAP_HOTPLUG_SURPRISE                => "FALSE",
      SLOT_CAP_MRL_SENSOR_PRESENT              => "FALSE",
      SLOT_CAP_NO_CMD_COMPLETED_SUPPORT        => "FALSE",
      SLOT_CAP_PHYSICAL_SLOT_NUM               => conv_integer(x"0000"),
      SLOT_CAP_POWER_CONTROLLER_PRESENT        => "FALSE",
      SLOT_CAP_POWER_INDICATOR_PRESENT         => "FALSE",
      SLOT_CAP_SLOT_POWER_LIMIT_SCALE          => 0,
      SLOT_CAP_SLOT_POWER_LIMIT_VALUE          => conv_integer(x"00"),
      TL_RX_RAM_RADDR_LATENCY                  => 0,
      TL_RX_RAM_RDATA_LATENCY                  => 2,
      TL_RX_RAM_WRITE_LATENCY                  => 0,
      TL_TX_RAM_RADDR_LATENCY                  => 0,
      TL_TX_RAM_RDATA_LATENCY                  => 2,
      TL_TX_RAM_WRITE_LATENCY                  => 0,

      UPCONFIG_CAPABLE                         => "TRUE",
      UPSTREAM_FACING                          => UPSTREAM_FACING,
      USER_CLK_FREQ                            => USER_CLK_FREQ,
      VC_BASE_PTR                              => conv_integer(x"10C"),
      VC_CAP_NEXTPTR                           => conv_integer(x"000"),
      VC_CAP_ON                                => "FALSE",
      VC_CAP_REJECT_SNOOP_TRANSACTIONS         => "FALSE",

      VC0_CPL_INFINITE                         => "TRUE",
      VC0_RX_RAM_LIMIT                         => VC0_RX_RAM_LIMIT,
      VC0_TOTAL_CREDITS_CD                     => VC0_TOTAL_CREDITS_CD,
      VC0_TOTAL_CREDITS_CH                     => VC0_TOTAL_CREDITS_CH,
      VC0_TOTAL_CREDITS_NPH                    => VC0_TOTAL_CREDITS_NPH,
      VC0_TOTAL_CREDITS_PD                     => VC0_TOTAL_CREDITS_PD,
      VC0_TOTAL_CREDITS_PH                     => 32,
      VC0_TX_LASTPACKET                        => 28,
      VENDOR_ID                                => conv_integer(C_VENDOR_ID),
      VSEC_BASE_PTR                            => conv_integer(x"000"),
      VSEC_CAP_NEXTPTR                         => conv_integer(x"000"),
      VSEC_CAP_ON                              => "FALSE",

      ALLOW_X8_GEN2                            => "FALSE",
      AER_BASE_PTR                             => conv_integer(x"000"),
      AER_CAP_ECRC_CHECK_CAPABLE               => "FALSE",
      AER_CAP_ECRC_GEN_CAPABLE                 => "FALSE",
      AER_CAP_ID                               => conv_integer(x"0001"),
      AER_CAP_INT_MSG_NUM_MSI                  => conv_integer(x"0a"),
      AER_CAP_INT_MSG_NUM_MSIX                 => conv_integer(x"15"),
      AER_CAP_NEXTPTR                          => conv_integer(x"160"),
      AER_CAP_ON                               => "FALSE",
      AER_CAP_PERMIT_ROOTERR_UPDATE            => "TRUE",
      AER_CAP_VERSION                          => conv_integer(x"1"),

      CAPABILITIES_PTR                         => conv_integer(x"40"),
      CRM_MODULE_RSTS                          => conv_integer(x"00"),
      DEV_CAP_ENDPOINT_L0S_LATENCY             => 0,
      DEV_CAP_ENDPOINT_L1_LATENCY              => 0,
      DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE     => "FALSE",
      DEV_CAP_ROLE_BASED_ERROR                 => "TRUE",
      DEV_CAP_RSVD_14_12                       => 0,
      DEV_CAP_RSVD_17_16                       => 0,
      DEV_CAP_RSVD_31_29                       => 0,
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE      => "TRUE",
      DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE      => "TRUE",
      DEV_CONTROL_AUX_POWER_SUPPORTED          => "FALSE",

      DISABLE_ASPM_L1_TIMER                    => "FALSE",
      DISABLE_BAR_FILTERING                    => "FALSE",
      DISABLE_ID_CHECK                         => "FALSE",
      DISABLE_RX_TC_FILTER                     => "FALSE",
      DNSTREAM_LINK_NUM                        => conv_integer(x"00"),

      DS_PORT_HOT_RST                          => "FALSE",  -- FALSE - for ROOT PORT(default), TRUE - for DOWNSTREAM PORT 
      DSN_CAP_ID                               => conv_integer(x"0003"),
      DSN_CAP_VERSION                          => conv_integer(x"1"),
      ENTER_RVRY_EI_L0                         => "TRUE",
      INFER_EI                                 => conv_integer(x"00"),
      IS_SWITCH                                => "FALSE",

      LAST_CONFIG_DWORD                        => conv_integer(x"042"),
      LINK_CAP_ASPM_SUPPORT                    => 1,
      LINK_CAP_CLOCK_POWER_MANAGEMENT          => "FALSE",
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1    => 7,
      LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2    => 7,
      LINK_CAP_L0S_EXIT_LATENCY_GEN1           => 7,
      LINK_CAP_L0S_EXIT_LATENCY_GEN2           => 7,
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1     => 7,
      LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2     => 7,
      LINK_CAP_L1_EXIT_LATENCY_GEN1            => 7,
      LINK_CAP_L1_EXIT_LATENCY_GEN2            => 7,
      LINK_CAP_RSVD_23_22                      => 0,

      MSI_BASE_PTR                             => conv_integer(x"48"),
      MSI_CAP_ID                               => conv_integer(x"05"),
      MSI_CAP_NEXTPTR                          => conv_integer(x"60"),
      MSIX_BASE_PTR                            => conv_integer(x"9c"),
      MSIX_CAP_ID                              => conv_integer(x"11"),
      MSIX_CAP_NEXTPTR                         => conv_integer(x"00"),
      N_FTS_COMCLK_GEN1                        => 255,
      N_FTS_COMCLK_GEN2                        => 254,
      N_FTS_GEN1                               => 255,
      N_FTS_GEN2                               => 255,

      PCIE_BASE_PTR                            => conv_integer(x"60"),
      PCIE_CAP_CAPABILITY_ID                   => conv_integer(x"10"),
      PCIE_CAP_CAPABILITY_VERSION              => PCIE_CAP_CAPABILITY_VERSION,
      PCIE_CAP_ON                              => "TRUE",
      PCIE_CAP_RSVD_15_14                      => 0,
      PCIE_CAP_SLOT_IMPLEMENTED                => CON_PCIE_CAP_SLOT_IMPLEMENTED,
      PCIE_REVISION                            => 2,
      PGL0_LANE                                => 0,
      PGL1_LANE                                => 1,
      PGL2_LANE                                => 2,
      PGL3_LANE                                => 3,
      PGL4_LANE                                => 4,
      PGL5_LANE                                => 5,
      PGL6_LANE                                => 6,
      PGL7_LANE                                => 7,
      PL_AUTO_CONFIG                           => 1,
      PL_FAST_TRAIN                            => C_PL_FAST_TRAIN_LOCAL,
      PCIE_EXT_CLK                             => PCIE_EXT_CLK,
      PCIE_EXT_GT_COMMON 		       => PCIE_EXT_GT_COMMON,
      EXT_CH_GT_DRP 			       => EXT_CH_GT_DRP,

      TX_MARGIN_FULL_0                         => conv_integer (x"4F"),
      TX_MARGIN_FULL_1                         => conv_integer (x"4e"),
      TX_MARGIN_FULL_2                         => conv_integer (x"4d"),
      TX_MARGIN_FULL_3                         => conv_integer (x"4c"),
      TX_MARGIN_FULL_4                         => conv_integer (x"43"),
      TX_MARGIN_LOW_0                          => conv_integer (x"45"),
      TX_MARGIN_LOW_1                          => conv_integer (x"46"),
      TX_MARGIN_LOW_2                          => conv_integer (x"43"),
      TX_MARGIN_LOW_3                          => conv_integer (x"42"),
      TX_MARGIN_LOW_4                          => conv_integer  (x"40"),
      PM_BASE_PTR                              => conv_integer(x"40"),
      PM_CAP_AUXCURRENT                        => 0,
      PM_CAP_ID                                => conv_integer(x"01"),
      PM_CAP_ON                                => "TRUE",
      PM_CAP_PME_CLOCK                         => "FALSE",
      PM_CAP_RSVD_04                           => 0,
      PM_CAP_VERSION                           => 3,
      PM_CSR_BPCCEN                            => "FALSE",
      PM_CSR_B2B3                              => "FALSE",
      RECRC_CHK                                => 0,
      RECRC_CHK_TRIM                           => "FALSE",
      SELECT_DLL_IF                            => "FALSE",
      SPARE_BIT1                               => 0,
      SPARE_BIT2                               => 0,
      SPARE_BIT3                               => 0,
      SPARE_BIT4                               => 0,
      SPARE_BIT5                               => 0,
      SPARE_BIT6                               => 0,
      SPARE_BIT7                               => 0,
      SPARE_BIT8                               => 0,
      SPARE_BYTE0                              => conv_integer(x"00"),
      SPARE_BYTE1                              => conv_integer(x"00"),
      SPARE_BYTE2                              => conv_integer(x"00"),
      SPARE_BYTE3                              => conv_integer(x"00"),
      SPARE_WORD0                              => conv_integer(x"00000000"),
      SPARE_WORD1                              => conv_integer(x"00000000"),
      SPARE_WORD2                              => conv_integer(x"00000000"),
      SPARE_WORD3                              => conv_integer(x"00000000"),

      TL_RBYPASS                               => "FALSE",
      TL_TFC_DISABLE                           => "FALSE",
      TL_TX_CHECKS_DISABLE                     => "FALSE",
      EXIT_LOOPBACK_ON_EI                      => "TRUE",
      UR_INV_REQ                               => "TRUE",

      VC_CAP_ID                                => conv_integer(x"0002"),
      VC_CAP_VERSION                           => conv_integer(x"1"),
      VSEC_CAP_HDR_ID                          => conv_integer(x"1234"),
      VSEC_CAP_HDR_LENGTH                      => conv_integer(x"018"),
      VSEC_CAP_HDR_REVISION                    => conv_integer(x"1"),
      VSEC_CAP_ID                              => conv_integer(x"000b"),
      VSEC_CAP_IS_LINK_VISIBLE                 => "FALSE",
      VSEC_CAP_VERSION                         => conv_integer(x"1"),
      C_BASEADDR_U                             => conv_integer(BASEADDR_U),-- AXI Lite Base Address upper
      C_BASEADDR_L                             => conv_integer(BASEADDR_L),-- AXI Lite Base Address lower
      C_HIGHADDR_U                             => conv_integer(HIGHADDR_U),-- AXI Lite High Address upper
      C_HIGHADDR_L                             => conv_integer(HIGHADDR_L),-- AXI Lite High Address lower
      C_MAX_LNK_WDT                            => 1,                    -- Maximum Number of PCIE Lanes
      C_ROOT_PORT                              => ROOT_PORT,            -- PCIe block is in root port mode
      C_RP_BAR_HIDE                            => C_RP_BAR_HIDE,        -- Hide RP PCIe BAR (prevent CPU from assigning address to RP BAR)
      C_RX_REALIGN                             => "FALSE",                -- Enable or Disable Realignment at RX Interface
      C_RX_PRESERVE_ORDER                      => "FALSE",               -- Preserve WR/ RD Ordering at the RX Interface
      C_LAST_CORE_CAP_ADDR                     => conv_integer(x"100"), -- DWORD address of last enabled block capability
      C_VSEC_CAP_ADDR                          => conv_integer(x"128"), -- DWORD address of start of VSEC Header
      C_VSEC_CAP_LAST                          => VSEC_CAP_LAST,
      C_VSEC_ID                                => conv_integer(x"0001"),
      C_DEVICE_NUMBER                          => 0,                    -- Device number for Root Port configurations only
      C_NUM_USER_INTR                          => NUM_OF_INTERRUPTS,
      C_USER_PTR                               => conv_integer(x"D8"),
      C_COMP_TIMEOUT                           => C_COMP_TIMEOUT,
      PTR_WIDTH                                => PTR_WIDTH,
      C_FAMILY                                 => FAMILY,
      USR_CFG                                  => "FALSE",
      USR_EXT_CFG                              => "FALSE",
      LINK_CAP_L0S_EXIT_LATENCY                => 7,
      LINK_CAP_L1_EXIT_LATENCY                 => 7,
      PLM_AUTO_CONFIG                          => "FALSE",
      FAST_TRAIN                               => C_PL_FAST_TRAIN_LOCAL,
      PCIE_GENERIC                             => PCIE_GENERIC, --conv_integer("000011101111"),
      GTP_SEL                                  => 0,
      CFG_VEN_ID                               => conv_integer(C_VENDOR_ID),
      CFG_DEV_ID                               => conv_integer(C_DEVICE_ID),
      CFG_REV_ID                               => conv_integer(C_REV_ID),
      CFG_SUBSYS_VEN_ID                        => conv_integer(C_SUBSYSTEM_VENDOR_ID),
      CFG_SUBSYS_ID                            => conv_integer(C_SUBSYSTEM_ID),

      AER_CAP_MULTIHEADER                      => "FALSE",
      AER_CAP_OPTIONAL_ERR_SUPPORT             => conv_integer(x"000000"),
      DEV_CAP2_ARI_FORWARDING_SUPPORTED        => "FALSE",
      DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED  => "FALSE",
      DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED  => "FALSE",
      DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED      => "FALSE",
      DEV_CAP2_CAS128_COMPLETER_SUPPORTED      => "FALSE",
      DEV_CAP2_TPH_COMPLETER_SUPPORTED         => conv_integer("00"),
      DEV_CONTROL_EXT_TAG_DEFAULT              => "FALSE",
      DISABLE_RX_POISONED_RESP                 => "FALSE",
      LINK_CAP_ASPM_OPTIONALITY                => "FALSE",
      RBAR_BASE_PTR                            => conv_integer(x"000"),
      RBAR_CAP_CONTROL_ENCODEDBAR0             => conv_integer(x"00"),
      RBAR_CAP_CONTROL_ENCODEDBAR1             => conv_integer(x"00"),
      RBAR_CAP_CONTROL_ENCODEDBAR2             => conv_integer(x"00"),
      RBAR_CAP_CONTROL_ENCODEDBAR3             => conv_integer(x"00"),
      RBAR_CAP_CONTROL_ENCODEDBAR4             => conv_integer(x"00"),
      RBAR_CAP_CONTROL_ENCODEDBAR5             => conv_integer(x"00"),
      RBAR_CAP_INDEX0                          => conv_integer(x"0"),
      RBAR_CAP_INDEX1                          => conv_integer(x"0"),
      RBAR_CAP_INDEX2                          => conv_integer(x"0"),
      RBAR_CAP_INDEX3                          => conv_integer(x"0"),
      RBAR_CAP_INDEX4                          => conv_integer(x"0"),
      RBAR_CAP_INDEX5                          => conv_integer(x"0"),
      RBAR_CAP_ON                              => "FALSE",
      RBAR_CAP_SUP0                            => conv_integer(x"00000001"),
      RBAR_CAP_SUP1                            => conv_integer(x"00000001"),
      RBAR_CAP_SUP2                            => conv_integer(x"00000001"),
      RBAR_CAP_SUP3                            => conv_integer(x"00000001"),
      RBAR_CAP_SUP4                            => conv_integer(x"00000001"),
      RBAR_CAP_SUP5                            => conv_integer(x"00000001"),
      RBAR_NUM                                 => conv_integer(x"0"),
      TRN_NP_FC                                => C_TRN_NP_FC, -- CR 824083
      TRN_DW                                   => TRN_DW,
      UR_ATOMIC                                => "FALSE",
      UR_PRS_RESPONSE                          => "TRUE",
      USER_CLK2_DIV2                           => USER_CLK2_DIV2,
      VC0_TOTAL_CREDITS_NPD                    => 24,
      LINK_CAP_RSVD_23                         => 0,
      CFG_ECRC_ERR_CPLSTAT                     => 0,
      DISABLE_ERR_MSG                          => "FALSE",
      DISABLE_LOCKED_FILTER                    => "FALSE",
      DISABLE_PPM_FILTER                       => "FALSE",
      ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED   => "FALSE",
      INTERRUPT_STAT_AUTO                      => "TRUE",
      MPS_FORCE                                => "FALSE",
      PM_ASPML0S_TIMEOUT                       => conv_integer(x"0000"),
      PM_ASPML0S_TIMEOUT_EN                    => "FALSE",
      PM_ASPML0S_TIMEOUT_FUNC                  => 0,
      PM_ASPM_FASTEXIT                         => "FALSE",
      PM_MF                                    => "FALSE",
      RP_AUTO_SPD                              => conv_integer(x"1"),
      RP_AUTO_SPD_LOOPCNT                      => conv_integer(x"1f"),
      SIM_VERSION                              => "1.0",
      SSL_MESSAGE_AUTO                         => "FALSE",
      TECRC_EP_INV                             => "FALSE",
      UR_CFG1                                  => "TRUE",
      USE_RID_PINS                             => "FALSE",
      DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED     => "FALSE",
      DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED    => "FALSE",
      DEV_CAP2_LTR_MECHANISM_SUPPORTED         => "FALSE",
      DEV_CAP2_MAX_ENDEND_TLP_PREFIXES         => conv_integer(x"0"),
      DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING      => "FALSE",
      RBAR_CAP_ID                              => conv_integer(x"0015"),
      RBAR_CAP_NEXTPTR                         => conv_integer(x"000"),
      RBAR_CAP_VERSION                         => conv_integer(x"1"),
      PCIE_USE_MODE                            => PCIE_USE_MODE,
      PCIE_GT_DEVICE                           => PCIE_GT_DEVICE,
      PCIE_CHAN_BOND                           => 0,
      PCIE_PLL_SEL                             => "CPLL",
      PCIE_ASYNC_EN                            => PCIE_ASYNC_EN,
      PCIE_TXBUF_EN                            => "FALSE"
      -- synthesis translate_off
      ,EXT_PIPE_INTERFACE                       =>  EXT_PIPE_INTERFACE
      -- synthesis translate_on
    )
    port map(
      -- 1. PCI Express (pci_exp) Interface
      ---------------------------------------------------------
      -- Tx
      pci_exp_txp                              => sig_pci_exp_txp,
      pci_exp_txn                              => sig_pci_exp_txn,
      -- Rx
      pci_exp_rxp                              => sig_pci_exp_rxp,
      pci_exp_rxn                              => sig_pci_exp_rxn,
qpll_drp_crscode      => qpll_drp_crscode    ,
  qpll_drp_fsm          => qpll_drp_fsm        ,
  qpll_drp_done         => qpll_drp_done       ,
  qpll_drp_reset        => qpll_drp_reset      ,
  qpll_qplllock         => qpll_qplllock       ,
  qpll_qplloutclk       => qpll_qplloutclk     ,
  qpll_qplloutrefclk    => qpll_qplloutrefclk  ,
   qpll_qplld    => qpll_qplld    ,
   qpll_qpllreset=> qpll_qpllreset,
   qpll_drp_clk  => qpll_drp_clk  ,
   qpll_drp_rst_n=> qpll_drp_rst_n,
   qpll_drp_ovrd => qpll_drp_ovrd ,
   qpll_drp_gen3 => qpll_drp_gen3 ,
   qpll_drp_start=> qpll_drp_start,

   pipe_txprbssel      => pipe_txprbssel     ,
   pipe_rxprbssel      => pipe_rxprbssel     ,
   pipe_txprbsforceerr => pipe_txprbsforceerr,
   pipe_rxprbscntreset => pipe_rxprbscntreset,
   pipe_loopback       => pipe_loopback      ,
   pipe_txinhibit        => pipe_txinhibit       ,

   pipe_rxprbserr        => pipe_rxprbserr       ,
   pipe_rst_fsm          => pipe_rst_fsm         ,
   pipe_qrst_fsm         => pipe_qrst_fsm        ,
   pipe_rate_fsm         => pipe_rate_fsm        ,
   pipe_sync_fsm_tx      => pipe_sync_fsm_tx     ,
   pipe_sync_fsm_rx      => pipe_sync_fsm_rx     ,
   pipe_drp_fsm          => pipe_drp_fsm         ,

   pipe_rst_idle => pipe_rst_idle ,
   pipe_qrst_idle=> pipe_qrst_idle,
   pipe_rate_idle=> pipe_rate_idle,
   pipe_eyescandataerror	=> pipe_eyescandataerror,
   pipe_rxstatus    => pipe_rxstatus,
   pipe_dmonitorout => pipe_dmonitorout,
  
   pipe_cpll_lock         =>  pipe_cpll_lock 	,
   pipe_qpll_lock         =>  pipe_qpll_lock 	,
   pipe_rxpmaresetdone    =>  pipe_rxpmaresetdone	,       
   pipe_rxbufstatus 	 =>  pipe_rxbufstatus 	,         
   pipe_txphaligndone     =>  pipe_txphaligndone 	,       
   pipe_txphinitdone 	 =>  pipe_txphinitdone 	,        
   pipe_txdlysresetdone   =>  pipe_txdlysresetdone,    
   pipe_rxphaligndone     =>  pipe_rxphaligndone 	,      
   pipe_rxdlysresetdone   =>  pipe_rxdlysresetdone,     
   pipe_rxsyncdone 	 =>  pipe_rxsyncdone 	,       
   pipe_rxdisperr 	 =>  pipe_rxdisperr 	,       
   pipe_rxnotintable 	 =>  pipe_rxnotintable 	,      
   pipe_rxcommadet 	 =>  pipe_rxcommadet 	,        

   gt_ch_drp_rdy => gt_ch_drp_rdy ,
   pipe_debug_0        => pipe_debug_0         ,
   pipe_debug_1        => pipe_debug_1         ,
   pipe_debug_2        => pipe_debug_2         ,
   pipe_debug_3        => pipe_debug_3         ,
   pipe_debug_4        => pipe_debug_4         ,
   pipe_debug_5        => pipe_debug_5         ,
   pipe_debug_6        => pipe_debug_6         ,
   pipe_debug_7        => pipe_debug_7         ,
   pipe_debug_8        => pipe_debug_8         ,
   pipe_debug_9        => pipe_debug_9         ,
   pipe_debug          => pipe_debug           ,

  common_commands_in		=>common_commands_in	,
  pipe_rx_0_sigs		=>pipe_rx_0_sigs	,
  pipe_rx_1_sigs		=>pipe_rx_1_sigs	,
  pipe_rx_2_sigs		=>pipe_rx_2_sigs	,
  pipe_rx_3_sigs		=>pipe_rx_3_sigs	,
  pipe_rx_4_sigs		=>pipe_rx_4_sigs	,
  pipe_rx_5_sigs		=>pipe_rx_5_sigs	,
  pipe_rx_6_sigs		=>pipe_rx_6_sigs	,
  pipe_rx_7_sigs		=>pipe_rx_7_sigs	,
                                                 
  common_commands_out		=>common_commands_out	,
  pipe_tx_0_sigs		=>pipe_tx_0_sigs	,
  pipe_tx_1_sigs		=>pipe_tx_1_sigs	,
  pipe_tx_2_sigs		=>pipe_tx_2_sigs	,
  pipe_tx_3_sigs		=>pipe_tx_3_sigs	,
  pipe_tx_4_sigs		=>pipe_tx_4_sigs	,
  pipe_tx_5_sigs		=>pipe_tx_5_sigs	,
  pipe_tx_6_sigs		=>pipe_tx_6_sigs	,
  pipe_tx_7_sigs		=>pipe_tx_7_sigs	,

INT_PCLK_OUT_SLAVE	=>		int_pclk_out_slave,	
INT_RXUSRCLK_OUT  	=>      	int_rxusrclk_out  ,      
INT_RXOUTCLK_OUT  	=>      	int_rxoutclk_out  ,      
INT_DCLK_OUT	  	=>      	int_dclk_out	  ,      
INT_USERCLK1_OUT  	=>      	int_userclk1_out  ,      
INT_USERCLK2_OUT  	=>      	int_userclk2_out  ,      
INT_OOBCLK_OUT	  	=>      	int_oobclk_out	  ,      
INT_MMCM_LOCK_OUT 	=>      	int_mmcm_lock_out ,      
INT_QPLLLOCK_OUT  	=>      	int_qplllock_out  ,      
INT_QPLLOUTCLK_OUT	=>		int_qplloutclk_out,	
INT_QPLLOUTREFCLK_OUT		=>	int_qplloutrefclk_out,	
INT_PCLK_SEL_SLAVE		=>	int_pclk_sel_slave   ,   

    -------------Channel DRP---------------------------------
   ext_ch_gt_drpclk    => ext_ch_gt_drpclk ,
   ext_ch_gt_drpaddr   => ext_ch_gt_drpaddr,
   ext_ch_gt_drpen     => ext_ch_gt_drpen  ,
   ext_ch_gt_drpdi     => ext_ch_gt_drpdi  ,
   ext_ch_gt_drpwe     => ext_ch_gt_drpwe  ,

   ext_ch_gt_drpdo     => ext_ch_gt_drpdo  ,
   ext_ch_gt_drprdy    => ext_ch_gt_drprdy ,

      clk_fab_refclk                           => clk_fab_refclk  ,
      clk_pclk                                 => clk_pclk        ,
      clk_rxusrclk                             => clk_rxusrclk    ,
      clk_dclk                                 => clk_dclk        ,
      clk_userclk1                             => clk_userclk1    ,
      clk_userclk2                             => clk_userclk2    ,
      clk_oobclk_in                            => clk_oobclk_in   ,
      clk_mmcm_lock                            => clk_mmcm_lock   ,
      clk_txoutclk                             => clk_txoutclk    ,
      clk_rxoutclk                             => clk_rxoutclk    ,
      clk_pclk_sel                             => clk_pclk_sel    ,
      clk_gen3                                 => clk_gen3        ,
      PIPE_MMCM_RST_N                          => pipe_mmcm_rst_n,


      ---------------------------------------------------------
      -- 2. Transaction (TRN) Interface
      ---------------------------------------------------------
      -- Rx
      rx_np_ok                                 => sig_rx_np_ok, --: in  std_logic;
      rx_np_req                                => sig_rx_np_req,--: in  std_logic;
      
      ---------------------------------------------
      -- AXI TX - RW Interface
      -----------
      s_axis_rw_tdata                          => sig_m_axis_rw_tdata,
      s_axis_rw_tvalid                         => sig_m_axis_rw_tvalid,
      s_axis_rw_tready                         => sig_m_axis_rw_tready,
      s_axis_rw_tstrb                          => sig_m_axis_rw_tstrb,
      s_axis_rw_tlast                          => sig_m_axis_rw_tlast,
      s_axis_rw_tuser                          => "0000",

      -- AXI TX - RR Interface
      -------------
      s_axis_rr_tdata                          => sig_m_axis_rr_tdata,
      s_axis_rr_tvalid                         => sig_m_axis_rr_tvalid,
      s_axis_rr_tready                         => sig_m_axis_rr_tready,
      s_axis_rr_tstrb                          => sig_m_axis_rr_tstrb,
      s_axis_rr_tlast                          => sig_m_axis_rr_tlast,
      s_axis_rr_tuser                          => "0000",

      -- AXI TX - CC Interface
      -------------
      s_axis_cc_tdata                          => sig_m_axis_cc_tdata,
      s_axis_cc_tvalid                         => sig_m_axis_cc_tvalid,
      s_axis_cc_tready                         => sig_m_axis_cc_tready,
      s_axis_cc_tstrb                          => sig_m_axis_cc_tstrb,
      s_axis_cc_tlast                          => sig_m_axis_cc_tlast,
      s_axis_cc_tuser                          => sig_m_axis_cc_tuser(3 downto 0),

      -- AXI RX - CW Interface
      -------------
      m_axis_cw_tdata                          => sig_s_axis_cw_tdata,
      m_axis_cw_tvalid                         => sig_s_axis_cw_tvalid,
      m_axis_cw_tready                         => sig_s_axis_cw_tready,
      m_axis_cw_tstrb                          => sig_s_axis_cw_tstrb,
      m_axis_cw_tlast                          => sig_s_axis_cw_tlast,
      m_axis_cw_tuser                          => sig_s_axis_cw_tuser,
 
      -- AXI RX - CR Interface
      -------------
      m_axis_cr_tdata                          => sig_s_axis_cr_tdata,
      m_axis_cr_tvalid                         => sig_s_axis_cr_tvalid,
      m_axis_cr_tready                         => sig_s_axis_cr_tready,
      m_axis_cr_tstrb                          => sig_s_axis_cr_tstrb,
      m_axis_cr_tlast                          => sig_s_axis_cr_tlast,
      m_axis_cr_tuser                          => sig_s_axis_cr_tuser,

      -- AXI RX - RC Interface
      -------------
      m_axis_rc_tdata                          => sig_s_axis_rc_tdata,
      m_axis_rc_tvalid                         => sig_s_axis_rc_tvalid,
      m_axis_rc_tready                         => sig_s_axis_rc_tready,
      m_axis_rc_tstrb                          => sig_s_axis_rc_tstrb,
      m_axis_rc_tlast                          => sig_s_axis_rc_tlast,
      --m_axis_rc_tuser                          => 

      -- AXI -Lite Interface - CFG Block
      ---------------------------
      s_axi_ctl_awaddr                         => s_axi_ctl_awaddr, -- AXI Lite Write address
      s_axi_ctl_awvalid                        => s_axi_ctl_awvalid,-- AXI Lite Write Address Valid
      s_axi_ctl_awready                        => s_axi_ctl_awready,-- AXI Lite Write Address Core ready
      s_axi_ctl_wdata                          => s_axi_ctl_wdata,  -- AXI Lite Write Data
      s_axi_ctl_wstrb                          => s_axi_ctl_wstrb,  -- AXI Lite Write Data strobe
      s_axi_ctl_wvalid                         => s_axi_ctl_wvalid, -- AXI Lite Write data Valid
      s_axi_ctl_wready                         => s_axi_ctl_wready, -- AXI Lite Write Data Core ready
      s_axi_ctl_bresp                          => s_axi_ctl_bresp,  -- AXI Lite Write Data strobe
      s_axi_ctl_bvalid                         => s_axi_ctl_bvalid, -- AXI Lite Write data Valid
      s_axi_ctl_bready                         => s_axi_ctl_bready, -- AXI Lite Write Data Core ready

      s_axi_ctl_araddr                         => s_axi_ctl_araddr, -- AXI Lite Read address
      s_axi_ctl_arvalid                        => s_axi_ctl_arvalid,-- AXI Lite Read Address Valid
      s_axi_ctl_arready                        => s_axi_ctl_arready,-- AXI Lite Read Address Core ready
      s_axi_ctl_rdata                          => s_axi_ctl_rdata,  -- AXI Lite Read Data
      s_axi_ctl_rresp                          => s_axi_ctl_rresp,  -- AXI Lite Read Data strobe
      s_axi_ctl_rvalid                         => s_axi_ctl_rvalid, -- AXI Lite Read data Valid
      s_axi_ctl_rready                         => s_axi_ctl_rready, -- AXI Lite Read Data Core ready

      -- AXI Lite User IPIC Signals
      -----------------------------
      Bus2IP_CS                                => sig_Bus2IP_CS,    -- Chip Select
      Bus2IP_BE                                => sig_Bus2IP_BE,    -- Byte Enable Vector
      Bus2IP_RNW                               => sig_Bus2IP_RNW,   -- Read Npt Write Qualifier
      Bus2IP_Addr                              => sig_Bus2IP_Addr,  -- Address Bus
      Bus2IP_Data                              => sig_Bus2IP_Data,  -- Write Data Bus
      IP2Bus_RdAck                             => sig_IP2Bus_RdAck, -- Read Acknowledgement
      IP2Bus_WrAck                             => sig_IP2Bus_WrAck, -- Write Acknowledgement
      IP2Bus_Data                              => sig_IP2Bus_Data,  -- Read Data Bus
      IP2Bus_Error                             => sig_IP2Bus_Error, -- Error Qualifier

      --Interrupts
      -------------------
      ctl_intr                                 => interrupt_out,    -- user interrupt
      ctl_user_intr                            => interrupt_vector,
  
      -- User Misc.
      -------------
      --user_turnoff_ok                          => in  std_logic;                                 -- Turnoff OK from user
      --user_tcfg_gnt                            => in  std_logic;                                 -- Send cfg OK from user

      np_cpl_pending                           => np_cpl_pending_qual,-- in  std_logic;
      RP_bridge_en                             => RP_bridge_en,

      ---------------------------------------------------------
      -- 3. Configuration (CFG) Interface
      ---------------------------------------------------------

      blk_err_cor                              => '0',--in  std_logic;
      blk_err_ur                               => '0',--in  std_logic;
      blk_err_ecrc                             => '0',--in  std_logic;
      blk_err_cpl_timeout                      => '0',--in  std_logic;
      blk_err_cpl_abort                        => '0',--in  std_logic;
      blk_err_cpl_unexpect                     => '0',--in  std_logic;
      blk_err_posted                           => '0',--in  std_logic;
      blk_err_locked                           => '0',--in  std_logic;
      blk_err_tlp_cpl_header                   => x"0000_0000_0000",--in  std_logic_vector(47 downto 0);
      --blk_err_cpl_rdy                          => out std_logic;
      blk_interrupt                            => sig_blk_interrupt,--in  std_logic;
      --blk_interrupt                            => '0',--in  std_logic;
      blk_interrupt_rdy                        => sig_blk_interrupt_rdy, --out std_logic;
      blk_interrupt_assert                     => sig_blk_interrupt_assert,--in  std_logic;
      blk_interrupt_di                         => sig_blk_interrupt_di,--in  std_logic_vector(7 downto 0);
      --cfg_interrupt_do                         => out std_logic_vector(7 downto 0);
      blk_interrupt_mmenable                   => MSI_Vector_Width,
      blk_interrupt_msienable                  => sig_blk_interrupt_msienable, -- out std_logic;
      --blk_interrupt_msixenable                 => out std_logic;
      --blk_interrupt_msixfm                     => out std_logic;
      blk_trn_pending                          => '0',--in  std_logic;
      cfg_pm_send_pme_to                       => '0',--in  std_logic;
      --blk_status                               => out std_logic_vector(15 downto 0);
      blk_command                              => sig_blk_command,
      --blk_dstatus                              => out std_logic_vector(15 downto 0);
      blk_dcommand                             => sig_blk_dcontrol,
      blk_lstatus                              => sig_blk_lstatus,
      --blk_lcommand                             => out std_logic_vector(15 downto 0);
      --blk_dcommand2                            => out std_logic_vector(15 downto 0);

      --blk_pcie_link_state                      => out std_logic_vector(2 downto 0);
      blk_dsn                                  => x"0000000000000000",--in  std_logic_vector(63 downto 0);
      --blk_pmcsr_pme_en                         => out std_logic;
      --blk_pmcsr_pme_status                     => out std_logic;
      --blk_pmcsr_powerstate                     => out std_logic_vector(1 downto 0);

      --cfg_msg_received                         => out std_logic;
      --blk_msg_data                             => out std_logic_vector(15 downto 0);
      --blk_msg_received_err_cor                 => out std_logic;
      --blk_msg_received_err_non_fatal           => out std_logic;
      --blk_msg_received_err_fatal               => out std_logic;
      --blk_msg_received_pme_to_ack              => out std_logic;
      --blk_msg_received_assert_inta             => out std_logic;
      --blk_msg_received_assert_intb             => out std_logic;
      --blk_msg_received_assert_intc             => out std_logic;
      --blk_msg_received_assert_intd             => out std_logic;
      --blk_msg_received_deassert_inta           => out std_logic;
      --blk_msg_received_deassert_intb           => out std_logic;
      --blk_msg_received_deassert_intc           => out std_logic;
      --blk_msg_received_deassert_intd           => out std_logic;

      blk_link_up                              => sig_blk_lnk_up,

      blk_ds_bus_number                        => x"00",--in  std_logic_vector(7 downto 0);
      blk_ds_device_number                     => "00000",--in  std_logic_vector(4 downto 0);

      -- Only for End point Cores
      --blk_to_turnoff                           => out  std_logic;
      blk_turnoff_ok                           => '0',--in std_logic;
      blk_pm_wake                              => '0',--in std_logic;

      blk_bus_number                           => sig_blk_bus_number,
      blk_device_number                        => sig_blk_device_number,
      blk_function_number                      => sig_blk_function_number,

      ---------------------------------------------------------
      -- 4. Physical Layer Control and Status (PL) Interface
      ---------------------------------------------------------

      --blk_pl_initial_link_width                => out std_logic_vector(2 downto 0);
      --blk_pl_lane_reversal_mode                => out std_logic_vector(1 downto 0);
      --blk_pl_link_gen2_capable                 => out std_logic;
      --blk_pl_link_partner_gen2_supported       => out std_logic;
      --blk_pl_link_upcfg_capable                => out std_logic;
      --blk_pl_ltssm_state                       => out std_logic_vector(5 downto 0);
      --blk_pl_sel_link_rate                     => out std_logic;
      --blk_pl_sel_link_width                    => out std_logic_vector(1 downto 0);
      blk_pl_upstream_prefer_deemph            => '0',--in  std_logic;
      --blk_pl_hot_rst                           => out std_logic;

      -- Flow Control
      --blk_fc_cpld                              => out std_logic_vector(11 downto 0);
      --blk_fc_cplh                              => out std_logic_vector(7 downto 0);
      --blk_fc_npd                               => out std_logic_vector(11 downto 0);
      --blk_fc_nph                               => out std_logic_vector(7 downto 0);
      --blk_fc_pd                                => out std_logic_vector(11 downto 0);
      --blk_fc_ph                                => out std_logic_vector(7 downto 0);
      blk_fc_sel                               => "100",--in  std_logic_vector(2 downto 0);

      -- Tx

      --blk_tbuf_av                              => out std_logic_vector(5 downto 0);
      --blk_tcfg_req                             => out std_logic;                                    
      blk_tcfg_gnt                             => '1',--in  std_logic;                               

      --tx_err_drop                              => --out std_logic;

      --S-6 Specific

      --cfg_do                                   => out std_logic_vector(31 downto 0);
      --cfg_rd_wr_done                           => out std_logic;                                
      cfg_dwaddr                               => "0000000000",--in  std_logic_vector(9 downto 0);
      cfg_rd_en                                => '0',--in  std_logic;                          

      ---------------------------------------------------------
      -- 5. System  (SYS) Interface
      ---------------------------------------------------------

      com_sysclk                               => REFCLK,
      com_sysrst                               => axi_areset,
      mmcm_lock                                => sig_mmcm_lock,
      com_iclk                                 => sig_axi_aclk_out,
      com_cclk                                 => sig_axi_ctl_aclk_out,
      config_gen_req				=> config_gen_req
      --com_corereset                            => out std_logic,
      
    );


end architecture;



